-- Pyramic_Array.vhd

-- Generated using ACDS version 16.0 211

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Pyramic_Array is
	port (
		audio_0_external_interface_BCLK                  : in    std_logic                     := '0';             --                  audio_0_external_interface.BCLK
		audio_0_external_interface_DACDAT                : out   std_logic;                                        --                                            .DACDAT
		audio_0_external_interface_DACLRCK               : in    std_logic                     := '0';             --                                            .DACLRCK
		audio_and_video_config_0_external_interface_SDAT : inout std_logic                     := '0';             -- audio_and_video_config_0_external_interface.SDAT
		audio_and_video_config_0_external_interface_SCLK : out   std_logic;                                        --                                            .SCLK
		clk_clk                                          : in    std_logic                     := '0';             --                                         clk.clk
		hps_0_ddr_mem_a                                  : out   std_logic_vector(14 downto 0);                    --                                   hps_0_ddr.mem_a
		hps_0_ddr_mem_ba                                 : out   std_logic_vector(2 downto 0);                     --                                            .mem_ba
		hps_0_ddr_mem_ck                                 : out   std_logic;                                        --                                            .mem_ck
		hps_0_ddr_mem_ck_n                               : out   std_logic;                                        --                                            .mem_ck_n
		hps_0_ddr_mem_cke                                : out   std_logic;                                        --                                            .mem_cke
		hps_0_ddr_mem_cs_n                               : out   std_logic;                                        --                                            .mem_cs_n
		hps_0_ddr_mem_ras_n                              : out   std_logic;                                        --                                            .mem_ras_n
		hps_0_ddr_mem_cas_n                              : out   std_logic;                                        --                                            .mem_cas_n
		hps_0_ddr_mem_we_n                               : out   std_logic;                                        --                                            .mem_we_n
		hps_0_ddr_mem_reset_n                            : out   std_logic;                                        --                                            .mem_reset_n
		hps_0_ddr_mem_dq                                 : inout std_logic_vector(31 downto 0) := (others => '0'); --                                            .mem_dq
		hps_0_ddr_mem_dqs                                : inout std_logic_vector(3 downto 0)  := (others => '0'); --                                            .mem_dqs
		hps_0_ddr_mem_dqs_n                              : inout std_logic_vector(3 downto 0)  := (others => '0'); --                                            .mem_dqs_n
		hps_0_ddr_mem_odt                                : out   std_logic;                                        --                                            .mem_odt
		hps_0_ddr_mem_dm                                 : out   std_logic_vector(3 downto 0);                     --                                            .mem_dm
		hps_0_ddr_oct_rzqin                              : in    std_logic                     := '0';             --                                            .oct_rzqin
		hps_0_io_hps_io_emac1_inst_TX_CLK                : out   std_logic;                                        --                                    hps_0_io.hps_io_emac1_inst_TX_CLK
		hps_0_io_hps_io_emac1_inst_TXD0                  : out   std_logic;                                        --                                            .hps_io_emac1_inst_TXD0
		hps_0_io_hps_io_emac1_inst_TXD1                  : out   std_logic;                                        --                                            .hps_io_emac1_inst_TXD1
		hps_0_io_hps_io_emac1_inst_TXD2                  : out   std_logic;                                        --                                            .hps_io_emac1_inst_TXD2
		hps_0_io_hps_io_emac1_inst_TXD3                  : out   std_logic;                                        --                                            .hps_io_emac1_inst_TXD3
		hps_0_io_hps_io_emac1_inst_RXD0                  : in    std_logic                     := '0';             --                                            .hps_io_emac1_inst_RXD0
		hps_0_io_hps_io_emac1_inst_MDIO                  : inout std_logic                     := '0';             --                                            .hps_io_emac1_inst_MDIO
		hps_0_io_hps_io_emac1_inst_MDC                   : out   std_logic;                                        --                                            .hps_io_emac1_inst_MDC
		hps_0_io_hps_io_emac1_inst_RX_CTL                : in    std_logic                     := '0';             --                                            .hps_io_emac1_inst_RX_CTL
		hps_0_io_hps_io_emac1_inst_TX_CTL                : out   std_logic;                                        --                                            .hps_io_emac1_inst_TX_CTL
		hps_0_io_hps_io_emac1_inst_RX_CLK                : in    std_logic                     := '0';             --                                            .hps_io_emac1_inst_RX_CLK
		hps_0_io_hps_io_emac1_inst_RXD1                  : in    std_logic                     := '0';             --                                            .hps_io_emac1_inst_RXD1
		hps_0_io_hps_io_emac1_inst_RXD2                  : in    std_logic                     := '0';             --                                            .hps_io_emac1_inst_RXD2
		hps_0_io_hps_io_emac1_inst_RXD3                  : in    std_logic                     := '0';             --                                            .hps_io_emac1_inst_RXD3
		hps_0_io_hps_io_sdio_inst_CMD                    : inout std_logic                     := '0';             --                                            .hps_io_sdio_inst_CMD
		hps_0_io_hps_io_sdio_inst_D0                     : inout std_logic                     := '0';             --                                            .hps_io_sdio_inst_D0
		hps_0_io_hps_io_sdio_inst_D1                     : inout std_logic                     := '0';             --                                            .hps_io_sdio_inst_D1
		hps_0_io_hps_io_sdio_inst_CLK                    : out   std_logic;                                        --                                            .hps_io_sdio_inst_CLK
		hps_0_io_hps_io_sdio_inst_D2                     : inout std_logic                     := '0';             --                                            .hps_io_sdio_inst_D2
		hps_0_io_hps_io_sdio_inst_D3                     : inout std_logic                     := '0';             --                                            .hps_io_sdio_inst_D3
		hps_0_io_hps_io_uart0_inst_RX                    : in    std_logic                     := '0';             --                                            .hps_io_uart0_inst_RX
		hps_0_io_hps_io_uart0_inst_TX                    : out   std_logic;                                        --                                            .hps_io_uart0_inst_TX
		hps_0_io_hps_io_gpio_inst_GPIO35                 : inout std_logic                     := '0';             --                                            .hps_io_gpio_inst_GPIO35
		hps_0_io_hps_io_gpio_inst_GPIO53                 : inout std_logic                     := '0';             --                                            .hps_io_gpio_inst_GPIO53
		hps_0_io_hps_io_gpio_inst_GPIO54                 : inout std_logic                     := '0';             --                                            .hps_io_gpio_inst_GPIO54
		output_switcher_0_source_select_new_signal       : in    std_logic                     := '0';             --             output_switcher_0_source_select.new_signal
		output_switcher_0_source_select_new_signal_1     : in    std_logic                     := '0';             --                                            .new_signal_1
		output_switcher_1_source_select_new_signal       : in    std_logic                     := '0';             --             output_switcher_1_source_select.new_signal
		output_switcher_1_source_select_new_signal_1     : in    std_logic                     := '0';             --                                            .new_signal_1
		pll_0_outclk3_audio_clk                          : out   std_logic;                                        --                         pll_0_outclk3_audio.clk
		pll_0_sdram_clk                                  : out   std_logic;                                        --                                 pll_0_sdram.clk
		reset_reset_n                                    : in    std_logic                     := '0';             --                                       reset.reset_n
		spi_system_0_spi_interface_convst0               : out   std_logic;                                        --                  spi_system_0_spi_interface.convst0
		spi_system_0_spi_interface_convst1               : out   std_logic;                                        --                                            .convst1
		spi_system_0_spi_interface_convst2               : out   std_logic;                                        --                                            .convst2
		spi_system_0_spi_interface_cs0_n                 : out   std_logic;                                        --                                            .cs0_n
		spi_system_0_spi_interface_cs1_n                 : out   std_logic;                                        --                                            .cs1_n
		spi_system_0_spi_interface_cs2_n                 : out   std_logic;                                        --                                            .cs2_n
		spi_system_0_spi_interface_miso_00               : in    std_logic                     := '0';             --                                            .miso_00
		spi_system_0_spi_interface_miso_01               : in    std_logic                     := '0';             --                                            .miso_01
		spi_system_0_spi_interface_miso_10               : in    std_logic                     := '0';             --                                            .miso_10
		spi_system_0_spi_interface_miso_11               : in    std_logic                     := '0';             --                                            .miso_11
		spi_system_0_spi_interface_miso_20               : in    std_logic                     := '0';             --                                            .miso_20
		spi_system_0_spi_interface_miso_21               : in    std_logic                     := '0';             --                                            .miso_21
		spi_system_0_spi_interface_reset0                : out   std_logic;                                        --                                            .reset0
		spi_system_0_spi_interface_reset1                : out   std_logic;                                        --                                            .reset1
		spi_system_0_spi_interface_reset2                : out   std_logic;                                        --                                            .reset2
		spi_system_0_spi_interface_sclk0                 : out   std_logic;                                        --                                            .sclk0
		spi_system_0_spi_interface_sclk1                 : out   std_logic;                                        --                                            .sclk1
		spi_system_0_spi_interface_sclk2                 : out   std_logic;                                        --                                            .sclk2
		spi_system_0_spi_interface_busy_or0              : in    std_logic                     := '0';             --                                            .busy_or0
		spi_system_0_spi_interface_busy_or1              : in    std_logic                     := '0';             --                                            .busy_or1
		spi_system_0_spi_interface_busy_or2              : in    std_logic                     := '0'              --                                            .busy_or2
	);
end entity Pyramic_Array;

architecture rtl of Pyramic_Array is
	component Beamformer_Adder is
		generic (
			DATA_WIDTH : natural := 32
		);
		port (
			clk         : in  std_logic                     := 'X';             -- clk
			reset_n     : in  std_logic                     := 'X';             -- reset_n
			Audio_Ready : in  std_logic                     := 'X';             -- ready
			Audio_Valid : out std_logic;                                        -- valid
			Audio_data  : out std_logic_vector(31 downto 0);                    -- data
			FIR_data    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			FIR_Valid   : in  std_logic                     := 'X';             -- valid
			FIR_Ready   : out std_logic;                                        -- ready
			FIR_sop     : in  std_logic                     := 'X';             -- startofpacket
			FIR_eop     : in  std_logic                     := 'X';             -- endofpacket
			FIR_channel : in  std_logic_vector(5 downto 0)  := (others => 'X')  -- channel
		);
	end component Beamformer_Adder;

	component Pyramic_Array_FIR_LEFT is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset_n            : in  std_logic                     := 'X';             -- reset_n
			ast_sink_data      : in  std_logic_vector(21 downto 0) := (others => 'X'); -- data
			ast_sink_valid     : in  std_logic                     := 'X';             -- valid
			ast_sink_error     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- error
			ast_sink_sop       : in  std_logic                     := 'X';             -- startofpacket
			ast_sink_eop       : in  std_logic                     := 'X';             -- endofpacket
			ast_source_data    : out std_logic_vector(31 downto 0);                    -- data
			ast_source_valid   : out std_logic;                                        -- valid
			ast_source_error   : out std_logic_vector(1 downto 0);                     -- error
			ast_source_sop     : out std_logic;                                        -- startofpacket
			ast_source_eop     : out std_logic;                                        -- endofpacket
			ast_source_channel : out std_logic_vector(5 downto 0)                      -- channel
		);
	end component Pyramic_Array_FIR_LEFT;

	component Output_Buffer_Driver is
		generic (
			SAMPLE_WIDTH : natural := 32
		);
		port (
			clk                           : in  std_logic                     := 'X';             -- clk
			reset_n                       : in  std_logic                     := 'X';             -- reset_n
			Use_Memory                    : in  std_logic                     := 'X';             -- new_signal
			Is_LeftRight                  : in  std_logic                     := 'X';             -- new_signal_1
			DMA_Addr                      : out std_logic_vector(31 downto 0);                    -- address
			DMA_ByteEnable                : out std_logic_vector(3 downto 0);                     -- byteenable
			DMA_Read                      : out std_logic;                                        -- read
			DMA_Data                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			DMA_Valid                     : in  std_logic                     := 'X';             -- readdatavalid
			DMA_WaitRequest               : in  std_logic                     := 'X';             -- waitrequest
			In_Avalon_Ready               : out std_logic;                                        -- ready
			In_Avalon_Valid               : in  std_logic                     := 'X';             -- valid
			In_Avalon_Data                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			avalon_streaming_source_ready : in  std_logic                     := 'X';             -- ready
			avalon_streaming_source_data  : out std_logic_vector(31 downto 0);                    -- data
			avalon_streaming_source_valid : out std_logic                                         -- valid
		);
	end component Output_Buffer_Driver;

	component SPI_System is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset_n            : in  std_logic                     := 'X';             -- reset_n
			AM_Addr            : out std_logic_vector(31 downto 0);                    -- address
			AM_BurstCount      : out std_logic_vector(2 downto 0);                     -- burstcount
			AM_ByteEnable      : out std_logic_vector(3 downto 0);                     -- byteenable
			AM_DataWrite       : out std_logic_vector(31 downto 0);                    -- writedata
			AM_WaitRequest     : in  std_logic                     := 'X';             -- waitrequest
			AM_Write           : out std_logic;                                        -- write
			AS_Write           : in  std_logic                     := 'X';             -- write
			AS_Read            : in  std_logic                     := 'X';             -- read
			AS_ReadData        : out std_logic_vector(31 downto 0);                    -- readdata
			AS_WriteData       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			AS_Addr            : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			CONVST0            : out std_logic;                                        -- convst0
			CONVST1            : out std_logic;                                        -- convst1
			CONVST2            : out std_logic;                                        -- convst2
			CS0_n              : out std_logic;                                        -- cs0_n
			CS1_n              : out std_logic;                                        -- cs1_n
			CS2_n              : out std_logic;                                        -- cs2_n
			MISO_00            : in  std_logic                     := 'X';             -- miso_00
			MISO_01            : in  std_logic                     := 'X';             -- miso_01
			MISO_10            : in  std_logic                     := 'X';             -- miso_10
			MISO_11            : in  std_logic                     := 'X';             -- miso_11
			MISO_20            : in  std_logic                     := 'X';             -- miso_20
			MISO_21            : in  std_logic                     := 'X';             -- miso_21
			Reset0             : out std_logic;                                        -- reset0
			Reset1             : out std_logic;                                        -- reset1
			Reset2             : out std_logic;                                        -- reset2
			SCLK0              : out std_logic;                                        -- sclk0
			SCLK1              : out std_logic;                                        -- sclk1
			SCLK2              : out std_logic;                                        -- sclk2
			busy_OR0           : in  std_logic                     := 'X';             -- busy_or0
			busy_OR1           : in  std_logic                     := 'X';             -- busy_or1
			busy_OR2           : in  std_logic                     := 'X';             -- busy_or2
			Source_Data_Left   : out std_logic_vector(21 downto 0);                    -- data
			Source_sop_Left    : out std_logic;                                        -- startofpacket
			Source_eop_Left    : out std_logic;                                        -- endofpacket
			Source_Valid_Left  : out std_logic;                                        -- valid
			Source_Ready_Left  : in  std_logic                     := 'X';             -- ready
			Source_Data_Right  : out std_logic_vector(21 downto 0);                    -- data
			Source_Ready_Right : in  std_logic                     := 'X';             -- ready
			Source_Valid_Right : out std_logic;                                        -- valid
			Source_eop_Right   : out std_logic;                                        -- endofpacket
			Source_sop_Right   : out std_logic                                         -- startofpacket
		);
	end component SPI_System;

	component Pyramic_Array_audio_and_video_config_0 is
		port (
			clk         : in    std_logic                     := 'X';             -- clk
			reset       : in    std_logic                     := 'X';             -- reset
			address     : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			byteenable  : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			read        : in    std_logic                     := 'X';             -- read
			write       : in    std_logic                     := 'X';             -- write
			writedata   : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata    : out   std_logic_vector(31 downto 0);                    -- readdata
			waitrequest : out   std_logic;                                        -- waitrequest
			I2C_SDAT    : inout std_logic                     := 'X';             -- export
			I2C_SCLK    : out   std_logic                                         -- export
		);
	end component Pyramic_Array_audio_and_video_config_0;

	component Pyramic_Array_audio_controller is
		port (
			clk                          : in  std_logic                     := 'X';             -- clk
			reset                        : in  std_logic                     := 'X';             -- reset
			from_adc_left_channel_ready  : in  std_logic                     := 'X';             -- ready
			from_adc_left_channel_data   : out std_logic_vector(31 downto 0);                    -- data
			from_adc_left_channel_valid  : out std_logic;                                        -- valid
			from_adc_right_channel_ready : in  std_logic                     := 'X';             -- ready
			from_adc_right_channel_data  : out std_logic_vector(31 downto 0);                    -- data
			from_adc_right_channel_valid : out std_logic;                                        -- valid
			to_dac_left_channel_data     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			to_dac_left_channel_valid    : in  std_logic                     := 'X';             -- valid
			to_dac_left_channel_ready    : out std_logic;                                        -- ready
			to_dac_right_channel_data    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			to_dac_right_channel_valid   : in  std_logic                     := 'X';             -- valid
			to_dac_right_channel_ready   : out std_logic;                                        -- ready
			AUD_BCLK                     : in  std_logic                     := 'X';             -- export
			AUD_DACDAT                   : out std_logic;                                        -- export
			AUD_DACLRCK                  : in  std_logic                     := 'X'              -- export
		);
	end component Pyramic_Array_audio_controller;

	component Pyramic_Array_hps_0 is
		generic (
			F2S_Width : integer := 2;
			S2F_Width : integer := 2
		);
		port (
			mem_a                    : out   std_logic_vector(14 downto 0);                    -- mem_a
			mem_ba                   : out   std_logic_vector(2 downto 0);                     -- mem_ba
			mem_ck                   : out   std_logic;                                        -- mem_ck
			mem_ck_n                 : out   std_logic;                                        -- mem_ck_n
			mem_cke                  : out   std_logic;                                        -- mem_cke
			mem_cs_n                 : out   std_logic;                                        -- mem_cs_n
			mem_ras_n                : out   std_logic;                                        -- mem_ras_n
			mem_cas_n                : out   std_logic;                                        -- mem_cas_n
			mem_we_n                 : out   std_logic;                                        -- mem_we_n
			mem_reset_n              : out   std_logic;                                        -- mem_reset_n
			mem_dq                   : inout std_logic_vector(31 downto 0) := (others => 'X'); -- mem_dq
			mem_dqs                  : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs
			mem_dqs_n                : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs_n
			mem_odt                  : out   std_logic;                                        -- mem_odt
			mem_dm                   : out   std_logic_vector(3 downto 0);                     -- mem_dm
			oct_rzqin                : in    std_logic                     := 'X';             -- oct_rzqin
			hps_io_emac1_inst_TX_CLK : out   std_logic;                                        -- hps_io_emac1_inst_TX_CLK
			hps_io_emac1_inst_TXD0   : out   std_logic;                                        -- hps_io_emac1_inst_TXD0
			hps_io_emac1_inst_TXD1   : out   std_logic;                                        -- hps_io_emac1_inst_TXD1
			hps_io_emac1_inst_TXD2   : out   std_logic;                                        -- hps_io_emac1_inst_TXD2
			hps_io_emac1_inst_TXD3   : out   std_logic;                                        -- hps_io_emac1_inst_TXD3
			hps_io_emac1_inst_RXD0   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD0
			hps_io_emac1_inst_MDIO   : inout std_logic                     := 'X';             -- hps_io_emac1_inst_MDIO
			hps_io_emac1_inst_MDC    : out   std_logic;                                        -- hps_io_emac1_inst_MDC
			hps_io_emac1_inst_RX_CTL : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RX_CTL
			hps_io_emac1_inst_TX_CTL : out   std_logic;                                        -- hps_io_emac1_inst_TX_CTL
			hps_io_emac1_inst_RX_CLK : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RX_CLK
			hps_io_emac1_inst_RXD1   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD1
			hps_io_emac1_inst_RXD2   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD2
			hps_io_emac1_inst_RXD3   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD3
			hps_io_sdio_inst_CMD     : inout std_logic                     := 'X';             -- hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK     : out   std_logic;                                        -- hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D3
			hps_io_uart0_inst_RX     : in    std_logic                     := 'X';             -- hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX     : out   std_logic;                                        -- hps_io_uart0_inst_TX
			hps_io_gpio_inst_GPIO35  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO35
			hps_io_gpio_inst_GPIO53  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO53
			hps_io_gpio_inst_GPIO54  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO54
			h2f_rst_n                : out   std_logic;                                        -- reset_n
			f2h_sdram0_clk           : in    std_logic                     := 'X';             -- clk
			f2h_sdram0_ADDRESS       : in    std_logic_vector(29 downto 0) := (others => 'X'); -- address
			f2h_sdram0_BURSTCOUNT    : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- burstcount
			f2h_sdram0_WAITREQUEST   : out   std_logic;                                        -- waitrequest
			f2h_sdram0_READDATA      : out   std_logic_vector(31 downto 0);                    -- readdata
			f2h_sdram0_READDATAVALID : out   std_logic;                                        -- readdatavalid
			f2h_sdram0_READ          : in    std_logic                     := 'X';             -- read
			f2h_sdram0_WRITEDATA     : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			f2h_sdram0_BYTEENABLE    : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			f2h_sdram0_WRITE         : in    std_logic                     := 'X';             -- write
			h2f_lw_axi_clk           : in    std_logic                     := 'X';             -- clk
			h2f_lw_AWID              : out   std_logic_vector(11 downto 0);                    -- awid
			h2f_lw_AWADDR            : out   std_logic_vector(20 downto 0);                    -- awaddr
			h2f_lw_AWLEN             : out   std_logic_vector(3 downto 0);                     -- awlen
			h2f_lw_AWSIZE            : out   std_logic_vector(2 downto 0);                     -- awsize
			h2f_lw_AWBURST           : out   std_logic_vector(1 downto 0);                     -- awburst
			h2f_lw_AWLOCK            : out   std_logic_vector(1 downto 0);                     -- awlock
			h2f_lw_AWCACHE           : out   std_logic_vector(3 downto 0);                     -- awcache
			h2f_lw_AWPROT            : out   std_logic_vector(2 downto 0);                     -- awprot
			h2f_lw_AWVALID           : out   std_logic;                                        -- awvalid
			h2f_lw_AWREADY           : in    std_logic                     := 'X';             -- awready
			h2f_lw_WID               : out   std_logic_vector(11 downto 0);                    -- wid
			h2f_lw_WDATA             : out   std_logic_vector(31 downto 0);                    -- wdata
			h2f_lw_WSTRB             : out   std_logic_vector(3 downto 0);                     -- wstrb
			h2f_lw_WLAST             : out   std_logic;                                        -- wlast
			h2f_lw_WVALID            : out   std_logic;                                        -- wvalid
			h2f_lw_WREADY            : in    std_logic                     := 'X';             -- wready
			h2f_lw_BID               : in    std_logic_vector(11 downto 0) := (others => 'X'); -- bid
			h2f_lw_BRESP             : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			h2f_lw_BVALID            : in    std_logic                     := 'X';             -- bvalid
			h2f_lw_BREADY            : out   std_logic;                                        -- bready
			h2f_lw_ARID              : out   std_logic_vector(11 downto 0);                    -- arid
			h2f_lw_ARADDR            : out   std_logic_vector(20 downto 0);                    -- araddr
			h2f_lw_ARLEN             : out   std_logic_vector(3 downto 0);                     -- arlen
			h2f_lw_ARSIZE            : out   std_logic_vector(2 downto 0);                     -- arsize
			h2f_lw_ARBURST           : out   std_logic_vector(1 downto 0);                     -- arburst
			h2f_lw_ARLOCK            : out   std_logic_vector(1 downto 0);                     -- arlock
			h2f_lw_ARCACHE           : out   std_logic_vector(3 downto 0);                     -- arcache
			h2f_lw_ARPROT            : out   std_logic_vector(2 downto 0);                     -- arprot
			h2f_lw_ARVALID           : out   std_logic;                                        -- arvalid
			h2f_lw_ARREADY           : in    std_logic                     := 'X';             -- arready
			h2f_lw_RID               : in    std_logic_vector(11 downto 0) := (others => 'X'); -- rid
			h2f_lw_RDATA             : in    std_logic_vector(31 downto 0) := (others => 'X'); -- rdata
			h2f_lw_RRESP             : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			h2f_lw_RLAST             : in    std_logic                     := 'X';             -- rlast
			h2f_lw_RVALID            : in    std_logic                     := 'X';             -- rvalid
			h2f_lw_RREADY            : out   std_logic                                         -- rready
		);
	end component Pyramic_Array_hps_0;

	component Pyramic_Array_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component Pyramic_Array_jtag_uart_0;

	component Pyramic_Array_pll_0 is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			outclk_1 : out std_logic;        -- clk
			outclk_2 : out std_logic;        -- clk
			outclk_3 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component Pyramic_Array_pll_0;

	component Pyramic_Array_pll_1 is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component Pyramic_Array_pll_1;

	component Pyramic_Array_sysid is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component Pyramic_Array_sysid;

	component Pyramic_Array_mm_interconnect_0 is
		port (
			pll_0_outclk0_clk                                                  : in  std_logic                     := 'X';             -- clk
			hps_0_f2h_sdram0_data_translator_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			Output_Switcher_0_reset_reset_bridge_in_reset_reset                : in  std_logic                     := 'X';             -- reset
			Output_Switcher_0_DMA_address                                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			Output_Switcher_0_DMA_waitrequest                                  : out std_logic;                                        -- waitrequest
			Output_Switcher_0_DMA_byteenable                                   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			Output_Switcher_0_DMA_read                                         : in  std_logic                     := 'X';             -- read
			Output_Switcher_0_DMA_readdata                                     : out std_logic_vector(31 downto 0);                    -- readdata
			Output_Switcher_0_DMA_readdatavalid                                : out std_logic;                                        -- readdatavalid
			Output_Switcher_1_DMA_address                                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			Output_Switcher_1_DMA_waitrequest                                  : out std_logic;                                        -- waitrequest
			Output_Switcher_1_DMA_byteenable                                   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			Output_Switcher_1_DMA_read                                         : in  std_logic                     := 'X';             -- read
			Output_Switcher_1_DMA_readdata                                     : out std_logic_vector(31 downto 0);                    -- readdata
			Output_Switcher_1_DMA_readdatavalid                                : out std_logic;                                        -- readdatavalid
			SPI_System_0_avalon_master_address                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			SPI_System_0_avalon_master_waitrequest                             : out std_logic;                                        -- waitrequest
			SPI_System_0_avalon_master_burstcount                              : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			SPI_System_0_avalon_master_byteenable                              : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			SPI_System_0_avalon_master_write                                   : in  std_logic                     := 'X';             -- write
			SPI_System_0_avalon_master_writedata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			hps_0_f2h_sdram0_data_address                                      : out std_logic_vector(29 downto 0);                    -- address
			hps_0_f2h_sdram0_data_write                                        : out std_logic;                                        -- write
			hps_0_f2h_sdram0_data_read                                         : out std_logic;                                        -- read
			hps_0_f2h_sdram0_data_readdata                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			hps_0_f2h_sdram0_data_writedata                                    : out std_logic_vector(31 downto 0);                    -- writedata
			hps_0_f2h_sdram0_data_burstcount                                   : out std_logic_vector(7 downto 0);                     -- burstcount
			hps_0_f2h_sdram0_data_byteenable                                   : out std_logic_vector(3 downto 0);                     -- byteenable
			hps_0_f2h_sdram0_data_readdatavalid                                : in  std_logic                     := 'X';             -- readdatavalid
			hps_0_f2h_sdram0_data_waitrequest                                  : in  std_logic                     := 'X'              -- waitrequest
		);
	end component Pyramic_Array_mm_interconnect_0;

	component Pyramic_Array_mm_interconnect_1 is
		port (
			hps_0_h2f_lw_axi_master_awid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- awid
			hps_0_h2f_lw_axi_master_awaddr                                      : in  std_logic_vector(20 downto 0) := (others => 'X'); -- awaddr
			hps_0_h2f_lw_axi_master_awlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awlen
			hps_0_h2f_lw_axi_master_awsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			hps_0_h2f_lw_axi_master_awburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			hps_0_h2f_lw_axi_master_awlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awlock
			hps_0_h2f_lw_axi_master_awcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awcache
			hps_0_h2f_lw_axi_master_awprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			hps_0_h2f_lw_axi_master_awvalid                                     : in  std_logic                     := 'X';             -- awvalid
			hps_0_h2f_lw_axi_master_awready                                     : out std_logic;                                        -- awready
			hps_0_h2f_lw_axi_master_wid                                         : in  std_logic_vector(11 downto 0) := (others => 'X'); -- wid
			hps_0_h2f_lw_axi_master_wdata                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wdata
			hps_0_h2f_lw_axi_master_wstrb                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- wstrb
			hps_0_h2f_lw_axi_master_wlast                                       : in  std_logic                     := 'X';             -- wlast
			hps_0_h2f_lw_axi_master_wvalid                                      : in  std_logic                     := 'X';             -- wvalid
			hps_0_h2f_lw_axi_master_wready                                      : out std_logic;                                        -- wready
			hps_0_h2f_lw_axi_master_bid                                         : out std_logic_vector(11 downto 0);                    -- bid
			hps_0_h2f_lw_axi_master_bresp                                       : out std_logic_vector(1 downto 0);                     -- bresp
			hps_0_h2f_lw_axi_master_bvalid                                      : out std_logic;                                        -- bvalid
			hps_0_h2f_lw_axi_master_bready                                      : in  std_logic                     := 'X';             -- bready
			hps_0_h2f_lw_axi_master_arid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- arid
			hps_0_h2f_lw_axi_master_araddr                                      : in  std_logic_vector(20 downto 0) := (others => 'X'); -- araddr
			hps_0_h2f_lw_axi_master_arlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arlen
			hps_0_h2f_lw_axi_master_arsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			hps_0_h2f_lw_axi_master_arburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			hps_0_h2f_lw_axi_master_arlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arlock
			hps_0_h2f_lw_axi_master_arcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arcache
			hps_0_h2f_lw_axi_master_arprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			hps_0_h2f_lw_axi_master_arvalid                                     : in  std_logic                     := 'X';             -- arvalid
			hps_0_h2f_lw_axi_master_arready                                     : out std_logic;                                        -- arready
			hps_0_h2f_lw_axi_master_rid                                         : out std_logic_vector(11 downto 0);                    -- rid
			hps_0_h2f_lw_axi_master_rdata                                       : out std_logic_vector(31 downto 0);                    -- rdata
			hps_0_h2f_lw_axi_master_rresp                                       : out std_logic_vector(1 downto 0);                     -- rresp
			hps_0_h2f_lw_axi_master_rlast                                       : out std_logic;                                        -- rlast
			hps_0_h2f_lw_axi_master_rvalid                                      : out std_logic;                                        -- rvalid
			hps_0_h2f_lw_axi_master_rready                                      : in  std_logic                     := 'X';             -- rready
			pll_0_outclk0_clk                                                   : in  std_logic                     := 'X';             -- clk
			audio_and_video_config_0_reset_reset_bridge_in_reset_reset          : in  std_logic                     := 'X';             -- reset
			hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			audio_and_video_config_0_avalon_av_config_slave_address             : out std_logic_vector(1 downto 0);                     -- address
			audio_and_video_config_0_avalon_av_config_slave_write               : out std_logic;                                        -- write
			audio_and_video_config_0_avalon_av_config_slave_read                : out std_logic;                                        -- read
			audio_and_video_config_0_avalon_av_config_slave_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			audio_and_video_config_0_avalon_av_config_slave_writedata           : out std_logic_vector(31 downto 0);                    -- writedata
			audio_and_video_config_0_avalon_av_config_slave_byteenable          : out std_logic_vector(3 downto 0);                     -- byteenable
			audio_and_video_config_0_avalon_av_config_slave_waitrequest         : in  std_logic                     := 'X';             -- waitrequest
			SPI_System_0_avalon_slave_address                                   : out std_logic_vector(2 downto 0);                     -- address
			SPI_System_0_avalon_slave_write                                     : out std_logic;                                        -- write
			SPI_System_0_avalon_slave_read                                      : out std_logic;                                        -- read
			SPI_System_0_avalon_slave_readdata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			SPI_System_0_avalon_slave_writedata                                 : out std_logic_vector(31 downto 0)                     -- writedata
		);
	end component Pyramic_Array_mm_interconnect_1;

	component Pyramic_Array_avalon_st_adapter is
		generic (
			inBitsPerSymbol : integer := 8;
			inUsePackets    : integer := 0;
			inDataWidth     : integer := 8;
			inChannelWidth  : integer := 3;
			inErrorWidth    : integer := 2;
			inUseEmptyPort  : integer := 0;
			inUseValid      : integer := 1;
			inUseReady      : integer := 1;
			inReadyLatency  : integer := 0;
			outDataWidth    : integer := 32;
			outChannelWidth : integer := 3;
			outErrorWidth   : integer := 2;
			outUseEmptyPort : integer := 0;
			outUseValid     : integer := 1;
			outUseReady     : integer := 1;
			outReadyLatency : integer := 0
		);
		port (
			in_clk_0_clk        : in  std_logic                     := 'X';             -- clk
			in_rst_0_reset      : in  std_logic                     := 'X';             -- reset
			in_0_data           : in  std_logic_vector(21 downto 0) := (others => 'X'); -- data
			in_0_valid          : in  std_logic                     := 'X';             -- valid
			in_0_ready          : out std_logic;                                        -- ready
			in_0_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_0_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_0_data          : out std_logic_vector(21 downto 0);                    -- data
			out_0_valid         : out std_logic;                                        -- valid
			out_0_startofpacket : out std_logic;                                        -- startofpacket
			out_0_endofpacket   : out std_logic;                                        -- endofpacket
			out_0_error         : out std_logic_vector(1 downto 0)                      -- error
		);
	end component Pyramic_Array_avalon_st_adapter;

	component Pyramic_Array_avalon_st_adapter_002 is
		generic (
			inBitsPerSymbol : integer := 8;
			inUsePackets    : integer := 0;
			inDataWidth     : integer := 8;
			inChannelWidth  : integer := 3;
			inErrorWidth    : integer := 2;
			inUseEmptyPort  : integer := 0;
			inUseValid      : integer := 1;
			inUseReady      : integer := 1;
			inReadyLatency  : integer := 0;
			outDataWidth    : integer := 32;
			outChannelWidth : integer := 3;
			outErrorWidth   : integer := 2;
			outUseEmptyPort : integer := 0;
			outUseValid     : integer := 1;
			outUseReady     : integer := 1;
			outReadyLatency : integer := 0
		);
		port (
			in_clk_0_clk        : in  std_logic                     := 'X';             -- clk
			in_rst_0_reset      : in  std_logic                     := 'X';             -- reset
			in_0_data           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			in_0_valid          : in  std_logic                     := 'X';             -- valid
			in_0_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_0_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			in_0_error          : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- error
			in_0_channel        : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- channel
			out_0_data          : out std_logic_vector(31 downto 0);                    -- data
			out_0_valid         : out std_logic;                                        -- valid
			out_0_ready         : in  std_logic                     := 'X';             -- ready
			out_0_startofpacket : out std_logic;                                        -- startofpacket
			out_0_endofpacket   : out std_logic;                                        -- endofpacket
			out_0_channel       : out std_logic_vector(5 downto 0)                      -- channel
		);
	end component Pyramic_Array_avalon_st_adapter_002;

	component pyramic_array_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component pyramic_array_rst_controller;

	component pyramic_array_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component pyramic_array_rst_controller_001;

	signal output_switcher_0_audio_streaming_source_valid                                : std_logic;                     -- Output_Switcher_0:avalon_streaming_source_valid -> audio_controller:to_dac_left_channel_valid
	signal output_switcher_0_audio_streaming_source_data                                 : std_logic_vector(31 downto 0); -- Output_Switcher_0:avalon_streaming_source_data -> audio_controller:to_dac_left_channel_data
	signal output_switcher_0_audio_streaming_source_ready                                : std_logic;                     -- audio_controller:to_dac_left_channel_ready -> Output_Switcher_0:avalon_streaming_source_ready
	signal output_switcher_1_audio_streaming_source_valid                                : std_logic;                     -- Output_Switcher_1:avalon_streaming_source_valid -> audio_controller:to_dac_right_channel_valid
	signal output_switcher_1_audio_streaming_source_data                                 : std_logic_vector(31 downto 0); -- Output_Switcher_1:avalon_streaming_source_data -> audio_controller:to_dac_right_channel_data
	signal output_switcher_1_audio_streaming_source_ready                                : std_logic;                     -- audio_controller:to_dac_right_channel_ready -> Output_Switcher_1:avalon_streaming_source_ready
	signal beamformer_left_source_beam_valid                                             : std_logic;                     -- Beamformer_LEFT:Audio_Valid -> Output_Switcher_0:In_Avalon_Valid
	signal beamformer_left_source_beam_data                                              : std_logic_vector(31 downto 0); -- Beamformer_LEFT:Audio_data -> Output_Switcher_0:In_Avalon_Data
	signal beamformer_left_source_beam_ready                                             : std_logic;                     -- Output_Switcher_0:In_Avalon_Ready -> Beamformer_LEFT:Audio_Ready
	signal beamformer_right_source_beam_valid                                            : std_logic;                     -- Beamformer_RIGHT:Audio_Valid -> Output_Switcher_1:In_Avalon_Valid
	signal beamformer_right_source_beam_data                                             : std_logic_vector(31 downto 0); -- Beamformer_RIGHT:Audio_data -> Output_Switcher_1:In_Avalon_Data
	signal beamformer_right_source_beam_ready                                            : std_logic;                     -- Output_Switcher_1:In_Avalon_Ready -> Beamformer_RIGHT:Audio_Ready
	signal pll_0_outclk0_clk                                                             : std_logic;                     -- pll_0:outclk_0 -> [Beamformer_LEFT:clk, Beamformer_RIGHT:clk, FIR_LEFT:clk, FIR_RIGHT:clk, Output_Switcher_0:clk, Output_Switcher_1:clk, SPI_System_0:clk, audio_and_video_config_0:clk, audio_controller:clk, avalon_st_adapter:in_clk_0_clk, avalon_st_adapter_001:in_clk_0_clk, avalon_st_adapter_002:in_clk_0_clk, avalon_st_adapter_003:in_clk_0_clk, hps_0:f2h_sdram0_clk, hps_0:h2f_lw_axi_clk, jtag_uart_0:clk, mm_interconnect_0:pll_0_outclk0_clk, mm_interconnect_1:pll_0_outclk0_clk, pll_1:refclk, rst_controller:clk, rst_controller_001:clk, rst_controller_003:clk, sysid:clock]
	signal output_switcher_0_dma_readdata                                                : std_logic_vector(31 downto 0); -- mm_interconnect_0:Output_Switcher_0_DMA_readdata -> Output_Switcher_0:DMA_Data
	signal output_switcher_0_dma_waitrequest                                             : std_logic;                     -- mm_interconnect_0:Output_Switcher_0_DMA_waitrequest -> Output_Switcher_0:DMA_WaitRequest
	signal output_switcher_0_dma_address                                                 : std_logic_vector(31 downto 0); -- Output_Switcher_0:DMA_Addr -> mm_interconnect_0:Output_Switcher_0_DMA_address
	signal output_switcher_0_dma_byteenable                                              : std_logic_vector(3 downto 0);  -- Output_Switcher_0:DMA_ByteEnable -> mm_interconnect_0:Output_Switcher_0_DMA_byteenable
	signal output_switcher_0_dma_read                                                    : std_logic;                     -- Output_Switcher_0:DMA_Read -> mm_interconnect_0:Output_Switcher_0_DMA_read
	signal output_switcher_0_dma_readdatavalid                                           : std_logic;                     -- mm_interconnect_0:Output_Switcher_0_DMA_readdatavalid -> Output_Switcher_0:DMA_Valid
	signal output_switcher_1_dma_readdata                                                : std_logic_vector(31 downto 0); -- mm_interconnect_0:Output_Switcher_1_DMA_readdata -> Output_Switcher_1:DMA_Data
	signal output_switcher_1_dma_waitrequest                                             : std_logic;                     -- mm_interconnect_0:Output_Switcher_1_DMA_waitrequest -> Output_Switcher_1:DMA_WaitRequest
	signal output_switcher_1_dma_address                                                 : std_logic_vector(31 downto 0); -- Output_Switcher_1:DMA_Addr -> mm_interconnect_0:Output_Switcher_1_DMA_address
	signal output_switcher_1_dma_byteenable                                              : std_logic_vector(3 downto 0);  -- Output_Switcher_1:DMA_ByteEnable -> mm_interconnect_0:Output_Switcher_1_DMA_byteenable
	signal output_switcher_1_dma_read                                                    : std_logic;                     -- Output_Switcher_1:DMA_Read -> mm_interconnect_0:Output_Switcher_1_DMA_read
	signal output_switcher_1_dma_readdatavalid                                           : std_logic;                     -- mm_interconnect_0:Output_Switcher_1_DMA_readdatavalid -> Output_Switcher_1:DMA_Valid
	signal spi_system_0_avalon_master_waitrequest                                        : std_logic;                     -- mm_interconnect_0:SPI_System_0_avalon_master_waitrequest -> SPI_System_0:AM_WaitRequest
	signal spi_system_0_avalon_master_address                                            : std_logic_vector(31 downto 0); -- SPI_System_0:AM_Addr -> mm_interconnect_0:SPI_System_0_avalon_master_address
	signal spi_system_0_avalon_master_byteenable                                         : std_logic_vector(3 downto 0);  -- SPI_System_0:AM_ByteEnable -> mm_interconnect_0:SPI_System_0_avalon_master_byteenable
	signal spi_system_0_avalon_master_writedata                                          : std_logic_vector(31 downto 0); -- SPI_System_0:AM_DataWrite -> mm_interconnect_0:SPI_System_0_avalon_master_writedata
	signal spi_system_0_avalon_master_write                                              : std_logic;                     -- SPI_System_0:AM_Write -> mm_interconnect_0:SPI_System_0_avalon_master_write
	signal spi_system_0_avalon_master_burstcount                                         : std_logic_vector(2 downto 0);  -- SPI_System_0:AM_BurstCount -> mm_interconnect_0:SPI_System_0_avalon_master_burstcount
	signal mm_interconnect_0_hps_0_f2h_sdram0_data_readdata                              : std_logic_vector(31 downto 0); -- hps_0:f2h_sdram0_READDATA -> mm_interconnect_0:hps_0_f2h_sdram0_data_readdata
	signal mm_interconnect_0_hps_0_f2h_sdram0_data_waitrequest                           : std_logic;                     -- hps_0:f2h_sdram0_WAITREQUEST -> mm_interconnect_0:hps_0_f2h_sdram0_data_waitrequest
	signal mm_interconnect_0_hps_0_f2h_sdram0_data_address                               : std_logic_vector(29 downto 0); -- mm_interconnect_0:hps_0_f2h_sdram0_data_address -> hps_0:f2h_sdram0_ADDRESS
	signal mm_interconnect_0_hps_0_f2h_sdram0_data_read                                  : std_logic;                     -- mm_interconnect_0:hps_0_f2h_sdram0_data_read -> hps_0:f2h_sdram0_READ
	signal mm_interconnect_0_hps_0_f2h_sdram0_data_byteenable                            : std_logic_vector(3 downto 0);  -- mm_interconnect_0:hps_0_f2h_sdram0_data_byteenable -> hps_0:f2h_sdram0_BYTEENABLE
	signal mm_interconnect_0_hps_0_f2h_sdram0_data_readdatavalid                         : std_logic;                     -- hps_0:f2h_sdram0_READDATAVALID -> mm_interconnect_0:hps_0_f2h_sdram0_data_readdatavalid
	signal mm_interconnect_0_hps_0_f2h_sdram0_data_write                                 : std_logic;                     -- mm_interconnect_0:hps_0_f2h_sdram0_data_write -> hps_0:f2h_sdram0_WRITE
	signal mm_interconnect_0_hps_0_f2h_sdram0_data_writedata                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:hps_0_f2h_sdram0_data_writedata -> hps_0:f2h_sdram0_WRITEDATA
	signal mm_interconnect_0_hps_0_f2h_sdram0_data_burstcount                            : std_logic_vector(7 downto 0);  -- mm_interconnect_0:hps_0_f2h_sdram0_data_burstcount -> hps_0:f2h_sdram0_BURSTCOUNT
	signal hps_0_h2f_lw_axi_master_awburst                                               : std_logic_vector(1 downto 0);  -- hps_0:h2f_lw_AWBURST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awburst
	signal hps_0_h2f_lw_axi_master_arlen                                                 : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_ARLEN -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arlen
	signal hps_0_h2f_lw_axi_master_wstrb                                                 : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_WSTRB -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wstrb
	signal hps_0_h2f_lw_axi_master_wready                                                : std_logic;                     -- mm_interconnect_1:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	signal hps_0_h2f_lw_axi_master_rid                                                   : std_logic_vector(11 downto 0); -- mm_interconnect_1:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	signal hps_0_h2f_lw_axi_master_rready                                                : std_logic;                     -- hps_0:h2f_lw_RREADY -> mm_interconnect_1:hps_0_h2f_lw_axi_master_rready
	signal hps_0_h2f_lw_axi_master_awlen                                                 : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_AWLEN -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awlen
	signal hps_0_h2f_lw_axi_master_wid                                                   : std_logic_vector(11 downto 0); -- hps_0:h2f_lw_WID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wid
	signal hps_0_h2f_lw_axi_master_arcache                                               : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_ARCACHE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arcache
	signal hps_0_h2f_lw_axi_master_wvalid                                                : std_logic;                     -- hps_0:h2f_lw_WVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wvalid
	signal hps_0_h2f_lw_axi_master_araddr                                                : std_logic_vector(20 downto 0); -- hps_0:h2f_lw_ARADDR -> mm_interconnect_1:hps_0_h2f_lw_axi_master_araddr
	signal hps_0_h2f_lw_axi_master_arprot                                                : std_logic_vector(2 downto 0);  -- hps_0:h2f_lw_ARPROT -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arprot
	signal hps_0_h2f_lw_axi_master_awprot                                                : std_logic_vector(2 downto 0);  -- hps_0:h2f_lw_AWPROT -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awprot
	signal hps_0_h2f_lw_axi_master_wdata                                                 : std_logic_vector(31 downto 0); -- hps_0:h2f_lw_WDATA -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wdata
	signal hps_0_h2f_lw_axi_master_arvalid                                               : std_logic;                     -- hps_0:h2f_lw_ARVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arvalid
	signal hps_0_h2f_lw_axi_master_awcache                                               : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_AWCACHE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awcache
	signal hps_0_h2f_lw_axi_master_arid                                                  : std_logic_vector(11 downto 0); -- hps_0:h2f_lw_ARID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arid
	signal hps_0_h2f_lw_axi_master_arlock                                                : std_logic_vector(1 downto 0);  -- hps_0:h2f_lw_ARLOCK -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arlock
	signal hps_0_h2f_lw_axi_master_awlock                                                : std_logic_vector(1 downto 0);  -- hps_0:h2f_lw_AWLOCK -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awlock
	signal hps_0_h2f_lw_axi_master_awaddr                                                : std_logic_vector(20 downto 0); -- hps_0:h2f_lw_AWADDR -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awaddr
	signal hps_0_h2f_lw_axi_master_bresp                                                 : std_logic_vector(1 downto 0);  -- mm_interconnect_1:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	signal hps_0_h2f_lw_axi_master_arready                                               : std_logic;                     -- mm_interconnect_1:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	signal hps_0_h2f_lw_axi_master_rdata                                                 : std_logic_vector(31 downto 0); -- mm_interconnect_1:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	signal hps_0_h2f_lw_axi_master_awready                                               : std_logic;                     -- mm_interconnect_1:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	signal hps_0_h2f_lw_axi_master_arburst                                               : std_logic_vector(1 downto 0);  -- hps_0:h2f_lw_ARBURST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arburst
	signal hps_0_h2f_lw_axi_master_arsize                                                : std_logic_vector(2 downto 0);  -- hps_0:h2f_lw_ARSIZE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arsize
	signal hps_0_h2f_lw_axi_master_bready                                                : std_logic;                     -- hps_0:h2f_lw_BREADY -> mm_interconnect_1:hps_0_h2f_lw_axi_master_bready
	signal hps_0_h2f_lw_axi_master_rlast                                                 : std_logic;                     -- mm_interconnect_1:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	signal hps_0_h2f_lw_axi_master_wlast                                                 : std_logic;                     -- hps_0:h2f_lw_WLAST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wlast
	signal hps_0_h2f_lw_axi_master_rresp                                                 : std_logic_vector(1 downto 0);  -- mm_interconnect_1:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	signal hps_0_h2f_lw_axi_master_awid                                                  : std_logic_vector(11 downto 0); -- hps_0:h2f_lw_AWID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awid
	signal hps_0_h2f_lw_axi_master_bid                                                   : std_logic_vector(11 downto 0); -- mm_interconnect_1:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	signal hps_0_h2f_lw_axi_master_bvalid                                                : std_logic;                     -- mm_interconnect_1:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	signal hps_0_h2f_lw_axi_master_awsize                                                : std_logic_vector(2 downto 0);  -- hps_0:h2f_lw_AWSIZE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awsize
	signal hps_0_h2f_lw_axi_master_awvalid                                               : std_logic;                     -- hps_0:h2f_lw_AWVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awvalid
	signal hps_0_h2f_lw_axi_master_rvalid                                                : std_logic;                     -- mm_interconnect_1:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	signal mm_interconnect_1_audio_and_video_config_0_avalon_av_config_slave_readdata    : std_logic_vector(31 downto 0); -- audio_and_video_config_0:readdata -> mm_interconnect_1:audio_and_video_config_0_avalon_av_config_slave_readdata
	signal mm_interconnect_1_audio_and_video_config_0_avalon_av_config_slave_waitrequest : std_logic;                     -- audio_and_video_config_0:waitrequest -> mm_interconnect_1:audio_and_video_config_0_avalon_av_config_slave_waitrequest
	signal mm_interconnect_1_audio_and_video_config_0_avalon_av_config_slave_address     : std_logic_vector(1 downto 0);  -- mm_interconnect_1:audio_and_video_config_0_avalon_av_config_slave_address -> audio_and_video_config_0:address
	signal mm_interconnect_1_audio_and_video_config_0_avalon_av_config_slave_read        : std_logic;                     -- mm_interconnect_1:audio_and_video_config_0_avalon_av_config_slave_read -> audio_and_video_config_0:read
	signal mm_interconnect_1_audio_and_video_config_0_avalon_av_config_slave_byteenable  : std_logic_vector(3 downto 0);  -- mm_interconnect_1:audio_and_video_config_0_avalon_av_config_slave_byteenable -> audio_and_video_config_0:byteenable
	signal mm_interconnect_1_audio_and_video_config_0_avalon_av_config_slave_write       : std_logic;                     -- mm_interconnect_1:audio_and_video_config_0_avalon_av_config_slave_write -> audio_and_video_config_0:write
	signal mm_interconnect_1_audio_and_video_config_0_avalon_av_config_slave_writedata   : std_logic_vector(31 downto 0); -- mm_interconnect_1:audio_and_video_config_0_avalon_av_config_slave_writedata -> audio_and_video_config_0:writedata
	signal mm_interconnect_1_spi_system_0_avalon_slave_readdata                          : std_logic_vector(31 downto 0); -- SPI_System_0:AS_ReadData -> mm_interconnect_1:SPI_System_0_avalon_slave_readdata
	signal mm_interconnect_1_spi_system_0_avalon_slave_address                           : std_logic_vector(2 downto 0);  -- mm_interconnect_1:SPI_System_0_avalon_slave_address -> SPI_System_0:AS_Addr
	signal mm_interconnect_1_spi_system_0_avalon_slave_read                              : std_logic;                     -- mm_interconnect_1:SPI_System_0_avalon_slave_read -> SPI_System_0:AS_Read
	signal mm_interconnect_1_spi_system_0_avalon_slave_write                             : std_logic;                     -- mm_interconnect_1:SPI_System_0_avalon_slave_write -> SPI_System_0:AS_Write
	signal mm_interconnect_1_spi_system_0_avalon_slave_writedata                         : std_logic_vector(31 downto 0); -- mm_interconnect_1:SPI_System_0_avalon_slave_writedata -> SPI_System_0:AS_WriteData
	signal spi_system_0_source_left_valid                                                : std_logic;                     -- SPI_System_0:Source_Valid_Left -> avalon_st_adapter:in_0_valid
	signal spi_system_0_source_left_data                                                 : std_logic_vector(21 downto 0); -- SPI_System_0:Source_Data_Left -> avalon_st_adapter:in_0_data
	signal spi_system_0_source_left_ready                                                : std_logic;                     -- avalon_st_adapter:in_0_ready -> SPI_System_0:Source_Ready_Left
	signal spi_system_0_source_left_startofpacket                                        : std_logic;                     -- SPI_System_0:Source_sop_Left -> avalon_st_adapter:in_0_startofpacket
	signal spi_system_0_source_left_endofpacket                                          : std_logic;                     -- SPI_System_0:Source_eop_Left -> avalon_st_adapter:in_0_endofpacket
	signal avalon_st_adapter_out_0_valid                                                 : std_logic;                     -- avalon_st_adapter:out_0_valid -> FIR_LEFT:ast_sink_valid
	signal avalon_st_adapter_out_0_data                                                  : std_logic_vector(21 downto 0); -- avalon_st_adapter:out_0_data -> FIR_LEFT:ast_sink_data
	signal avalon_st_adapter_out_0_startofpacket                                         : std_logic;                     -- avalon_st_adapter:out_0_startofpacket -> FIR_LEFT:ast_sink_sop
	signal avalon_st_adapter_out_0_endofpacket                                           : std_logic;                     -- avalon_st_adapter:out_0_endofpacket -> FIR_LEFT:ast_sink_eop
	signal avalon_st_adapter_out_0_error                                                 : std_logic_vector(1 downto 0);  -- avalon_st_adapter:out_0_error -> FIR_LEFT:ast_sink_error
	signal spi_system_0_source_right_valid                                               : std_logic;                     -- SPI_System_0:Source_Valid_Right -> avalon_st_adapter_001:in_0_valid
	signal spi_system_0_source_right_data                                                : std_logic_vector(21 downto 0); -- SPI_System_0:Source_Data_Right -> avalon_st_adapter_001:in_0_data
	signal spi_system_0_source_right_ready                                               : std_logic;                     -- avalon_st_adapter_001:in_0_ready -> SPI_System_0:Source_Ready_Right
	signal spi_system_0_source_right_startofpacket                                       : std_logic;                     -- SPI_System_0:Source_sop_Right -> avalon_st_adapter_001:in_0_startofpacket
	signal spi_system_0_source_right_endofpacket                                         : std_logic;                     -- SPI_System_0:Source_eop_Right -> avalon_st_adapter_001:in_0_endofpacket
	signal avalon_st_adapter_001_out_0_valid                                             : std_logic;                     -- avalon_st_adapter_001:out_0_valid -> FIR_RIGHT:ast_sink_valid
	signal avalon_st_adapter_001_out_0_data                                              : std_logic_vector(21 downto 0); -- avalon_st_adapter_001:out_0_data -> FIR_RIGHT:ast_sink_data
	signal avalon_st_adapter_001_out_0_startofpacket                                     : std_logic;                     -- avalon_st_adapter_001:out_0_startofpacket -> FIR_RIGHT:ast_sink_sop
	signal avalon_st_adapter_001_out_0_endofpacket                                       : std_logic;                     -- avalon_st_adapter_001:out_0_endofpacket -> FIR_RIGHT:ast_sink_eop
	signal avalon_st_adapter_001_out_0_error                                             : std_logic_vector(1 downto 0);  -- avalon_st_adapter_001:out_0_error -> FIR_RIGHT:ast_sink_error
	signal fir_left_avalon_streaming_source_valid                                        : std_logic;                     -- FIR_LEFT:ast_source_valid -> avalon_st_adapter_002:in_0_valid
	signal fir_left_avalon_streaming_source_data                                         : std_logic_vector(31 downto 0); -- FIR_LEFT:ast_source_data -> avalon_st_adapter_002:in_0_data
	signal fir_left_avalon_streaming_source_channel                                      : std_logic_vector(5 downto 0);  -- FIR_LEFT:ast_source_channel -> avalon_st_adapter_002:in_0_channel
	signal fir_left_avalon_streaming_source_startofpacket                                : std_logic;                     -- FIR_LEFT:ast_source_sop -> avalon_st_adapter_002:in_0_startofpacket
	signal fir_left_avalon_streaming_source_error                                        : std_logic_vector(1 downto 0);  -- FIR_LEFT:ast_source_error -> avalon_st_adapter_002:in_0_error
	signal fir_left_avalon_streaming_source_endofpacket                                  : std_logic;                     -- FIR_LEFT:ast_source_eop -> avalon_st_adapter_002:in_0_endofpacket
	signal avalon_st_adapter_002_out_0_valid                                             : std_logic;                     -- avalon_st_adapter_002:out_0_valid -> Beamformer_LEFT:FIR_Valid
	signal avalon_st_adapter_002_out_0_data                                              : std_logic_vector(31 downto 0); -- avalon_st_adapter_002:out_0_data -> Beamformer_LEFT:FIR_data
	signal avalon_st_adapter_002_out_0_ready                                             : std_logic;                     -- Beamformer_LEFT:FIR_Ready -> avalon_st_adapter_002:out_0_ready
	signal avalon_st_adapter_002_out_0_channel                                           : std_logic_vector(5 downto 0);  -- avalon_st_adapter_002:out_0_channel -> Beamformer_LEFT:FIR_channel
	signal avalon_st_adapter_002_out_0_startofpacket                                     : std_logic;                     -- avalon_st_adapter_002:out_0_startofpacket -> Beamformer_LEFT:FIR_sop
	signal avalon_st_adapter_002_out_0_endofpacket                                       : std_logic;                     -- avalon_st_adapter_002:out_0_endofpacket -> Beamformer_LEFT:FIR_eop
	signal fir_right_avalon_streaming_source_valid                                       : std_logic;                     -- FIR_RIGHT:ast_source_valid -> avalon_st_adapter_003:in_0_valid
	signal fir_right_avalon_streaming_source_data                                        : std_logic_vector(31 downto 0); -- FIR_RIGHT:ast_source_data -> avalon_st_adapter_003:in_0_data
	signal fir_right_avalon_streaming_source_channel                                     : std_logic_vector(5 downto 0);  -- FIR_RIGHT:ast_source_channel -> avalon_st_adapter_003:in_0_channel
	signal fir_right_avalon_streaming_source_startofpacket                               : std_logic;                     -- FIR_RIGHT:ast_source_sop -> avalon_st_adapter_003:in_0_startofpacket
	signal fir_right_avalon_streaming_source_error                                       : std_logic_vector(1 downto 0);  -- FIR_RIGHT:ast_source_error -> avalon_st_adapter_003:in_0_error
	signal fir_right_avalon_streaming_source_endofpacket                                 : std_logic;                     -- FIR_RIGHT:ast_source_eop -> avalon_st_adapter_003:in_0_endofpacket
	signal avalon_st_adapter_003_out_0_valid                                             : std_logic;                     -- avalon_st_adapter_003:out_0_valid -> Beamformer_RIGHT:FIR_Valid
	signal avalon_st_adapter_003_out_0_data                                              : std_logic_vector(31 downto 0); -- avalon_st_adapter_003:out_0_data -> Beamformer_RIGHT:FIR_data
	signal avalon_st_adapter_003_out_0_ready                                             : std_logic;                     -- Beamformer_RIGHT:FIR_Ready -> avalon_st_adapter_003:out_0_ready
	signal avalon_st_adapter_003_out_0_channel                                           : std_logic_vector(5 downto 0);  -- avalon_st_adapter_003:out_0_channel -> Beamformer_RIGHT:FIR_channel
	signal avalon_st_adapter_003_out_0_startofpacket                                     : std_logic;                     -- avalon_st_adapter_003:out_0_startofpacket -> Beamformer_RIGHT:FIR_sop
	signal avalon_st_adapter_003_out_0_endofpacket                                       : std_logic;                     -- avalon_st_adapter_003:out_0_endofpacket -> Beamformer_RIGHT:FIR_eop
	signal rst_controller_reset_out_reset                                                : std_logic;                     -- rst_controller:reset_out -> [audio_and_video_config_0:reset, audio_controller:reset, avalon_st_adapter:in_rst_0_reset, avalon_st_adapter_001:in_rst_0_reset, avalon_st_adapter_002:in_rst_0_reset, avalon_st_adapter_003:in_rst_0_reset, mm_interconnect_0:Output_Switcher_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:audio_and_video_config_0_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in]
	signal rst_controller_001_reset_out_reset                                            : std_logic;                     -- rst_controller_001:reset_out -> rst_controller_001_reset_out_reset:in
	signal hps_0_h2f_reset_reset                                                         : std_logic;                     -- hps_0:h2f_rst_n -> hps_0_h2f_reset_reset:in
	signal rst_controller_002_reset_out_reset                                            : std_logic;                     -- rst_controller_002:reset_out -> pll_0:rst
	signal rst_controller_003_reset_out_reset                                            : std_logic;                     -- rst_controller_003:reset_out -> [mm_interconnect_0:hps_0_f2h_sdram0_data_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_1:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset]
	signal reset_reset_n_ports_inv                                                       : std_logic;                     -- reset_reset_n:inv -> [pll_1:rst, rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0]
	signal rst_controller_reset_out_reset_ports_inv                                      : std_logic;                     -- rst_controller_reset_out_reset:inv -> [Beamformer_LEFT:reset_n, Beamformer_RIGHT:reset_n, FIR_LEFT:reset_n, FIR_RIGHT:reset_n, Output_Switcher_0:reset_n, Output_Switcher_1:reset_n, SPI_System_0:reset_n]
	signal rst_controller_001_reset_out_reset_ports_inv                                  : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> [jtag_uart_0:rst_n, sysid:reset_n]
	signal hps_0_h2f_reset_reset_ports_inv                                               : std_logic;                     -- hps_0_h2f_reset_reset:inv -> [rst_controller_001:reset_in1, rst_controller_002:reset_in1, rst_controller_003:reset_in0]

begin

	beamformer_left : component Beamformer_Adder
		generic map (
			DATA_WIDTH => 32
		)
		port map (
			clk         => pll_0_outclk0_clk,                         --       clock.clk
			reset_n     => rst_controller_reset_out_reset_ports_inv,  --       reset.reset_n
			Audio_Ready => beamformer_left_source_beam_ready,         -- Source_Beam.ready
			Audio_Valid => beamformer_left_source_beam_valid,         --            .valid
			Audio_data  => beamformer_left_source_beam_data,          --            .data
			FIR_data    => avalon_st_adapter_002_out_0_data,          --    Sink_FIR.data
			FIR_Valid   => avalon_st_adapter_002_out_0_valid,         --            .valid
			FIR_Ready   => avalon_st_adapter_002_out_0_ready,         --            .ready
			FIR_sop     => avalon_st_adapter_002_out_0_startofpacket, --            .startofpacket
			FIR_eop     => avalon_st_adapter_002_out_0_endofpacket,   --            .endofpacket
			FIR_channel => avalon_st_adapter_002_out_0_channel        --            .channel
		);

	beamformer_right : component Beamformer_Adder
		generic map (
			DATA_WIDTH => 32
		)
		port map (
			clk         => pll_0_outclk0_clk,                         --       clock.clk
			reset_n     => rst_controller_reset_out_reset_ports_inv,  --       reset.reset_n
			Audio_Ready => beamformer_right_source_beam_ready,        -- Source_Beam.ready
			Audio_Valid => beamformer_right_source_beam_valid,        --            .valid
			Audio_data  => beamformer_right_source_beam_data,         --            .data
			FIR_data    => avalon_st_adapter_003_out_0_data,          --    Sink_FIR.data
			FIR_Valid   => avalon_st_adapter_003_out_0_valid,         --            .valid
			FIR_Ready   => avalon_st_adapter_003_out_0_ready,         --            .ready
			FIR_sop     => avalon_st_adapter_003_out_0_startofpacket, --            .startofpacket
			FIR_eop     => avalon_st_adapter_003_out_0_endofpacket,   --            .endofpacket
			FIR_channel => avalon_st_adapter_003_out_0_channel        --            .channel
		);

	fir_left : component Pyramic_Array_FIR_LEFT
		port map (
			clk                => pll_0_outclk0_clk,                              --                     clk.clk
			reset_n            => rst_controller_reset_out_reset_ports_inv,       --                     rst.reset_n
			ast_sink_data      => avalon_st_adapter_out_0_data,                   --   avalon_streaming_sink.data
			ast_sink_valid     => avalon_st_adapter_out_0_valid,                  --                        .valid
			ast_sink_error     => avalon_st_adapter_out_0_error,                  --                        .error
			ast_sink_sop       => avalon_st_adapter_out_0_startofpacket,          --                        .startofpacket
			ast_sink_eop       => avalon_st_adapter_out_0_endofpacket,            --                        .endofpacket
			ast_source_data    => fir_left_avalon_streaming_source_data,          -- avalon_streaming_source.data
			ast_source_valid   => fir_left_avalon_streaming_source_valid,         --                        .valid
			ast_source_error   => fir_left_avalon_streaming_source_error,         --                        .error
			ast_source_sop     => fir_left_avalon_streaming_source_startofpacket, --                        .startofpacket
			ast_source_eop     => fir_left_avalon_streaming_source_endofpacket,   --                        .endofpacket
			ast_source_channel => fir_left_avalon_streaming_source_channel        --                        .channel
		);

	fir_right : component Pyramic_Array_FIR_LEFT
		port map (
			clk                => pll_0_outclk0_clk,                               --                     clk.clk
			reset_n            => rst_controller_reset_out_reset_ports_inv,        --                     rst.reset_n
			ast_sink_data      => avalon_st_adapter_001_out_0_data,                --   avalon_streaming_sink.data
			ast_sink_valid     => avalon_st_adapter_001_out_0_valid,               --                        .valid
			ast_sink_error     => avalon_st_adapter_001_out_0_error,               --                        .error
			ast_sink_sop       => avalon_st_adapter_001_out_0_startofpacket,       --                        .startofpacket
			ast_sink_eop       => avalon_st_adapter_001_out_0_endofpacket,         --                        .endofpacket
			ast_source_data    => fir_right_avalon_streaming_source_data,          -- avalon_streaming_source.data
			ast_source_valid   => fir_right_avalon_streaming_source_valid,         --                        .valid
			ast_source_error   => fir_right_avalon_streaming_source_error,         --                        .error
			ast_source_sop     => fir_right_avalon_streaming_source_startofpacket, --                        .startofpacket
			ast_source_eop     => fir_right_avalon_streaming_source_endofpacket,   --                        .endofpacket
			ast_source_channel => fir_right_avalon_streaming_source_channel        --                        .channel
		);

	output_switcher_0 : component Output_Buffer_Driver
		generic map (
			SAMPLE_WIDTH => 32
		)
		port map (
			clk                           => pll_0_outclk0_clk,                              --                  clock.clk
			reset_n                       => rst_controller_reset_out_reset_ports_inv,       --                  reset.reset_n
			Use_Memory                    => output_switcher_0_source_select_new_signal,     --          source_select.new_signal
			Is_LeftRight                  => output_switcher_0_source_select_new_signal_1,   --                       .new_signal_1
			DMA_Addr                      => output_switcher_0_dma_address,                  --                    DMA.address
			DMA_ByteEnable                => output_switcher_0_dma_byteenable,               --                       .byteenable
			DMA_Read                      => output_switcher_0_dma_read,                     --                       .read
			DMA_Data                      => output_switcher_0_dma_readdata,                 --                       .readdata
			DMA_Valid                     => output_switcher_0_dma_readdatavalid,            --                       .readdatavalid
			DMA_WaitRequest               => output_switcher_0_dma_waitrequest,              --                       .waitrequest
			In_Avalon_Ready               => beamformer_left_source_beam_ready,              --   Audio_Streaming_Sink.ready
			In_Avalon_Valid               => beamformer_left_source_beam_valid,              --                       .valid
			In_Avalon_Data                => beamformer_left_source_beam_data,               --                       .data
			avalon_streaming_source_ready => output_switcher_0_audio_streaming_source_ready, -- Audio_Streaming_Source.ready
			avalon_streaming_source_data  => output_switcher_0_audio_streaming_source_data,  --                       .data
			avalon_streaming_source_valid => output_switcher_0_audio_streaming_source_valid  --                       .valid
		);

	output_switcher_1 : component Output_Buffer_Driver
		generic map (
			SAMPLE_WIDTH => 32
		)
		port map (
			clk                           => pll_0_outclk0_clk,                              --                  clock.clk
			reset_n                       => rst_controller_reset_out_reset_ports_inv,       --                  reset.reset_n
			Use_Memory                    => output_switcher_1_source_select_new_signal,     --          source_select.new_signal
			Is_LeftRight                  => output_switcher_1_source_select_new_signal_1,   --                       .new_signal_1
			DMA_Addr                      => output_switcher_1_dma_address,                  --                    DMA.address
			DMA_ByteEnable                => output_switcher_1_dma_byteenable,               --                       .byteenable
			DMA_Read                      => output_switcher_1_dma_read,                     --                       .read
			DMA_Data                      => output_switcher_1_dma_readdata,                 --                       .readdata
			DMA_Valid                     => output_switcher_1_dma_readdatavalid,            --                       .readdatavalid
			DMA_WaitRequest               => output_switcher_1_dma_waitrequest,              --                       .waitrequest
			In_Avalon_Ready               => beamformer_right_source_beam_ready,             --   Audio_Streaming_Sink.ready
			In_Avalon_Valid               => beamformer_right_source_beam_valid,             --                       .valid
			In_Avalon_Data                => beamformer_right_source_beam_data,              --                       .data
			avalon_streaming_source_ready => output_switcher_1_audio_streaming_source_ready, -- Audio_Streaming_Source.ready
			avalon_streaming_source_data  => output_switcher_1_audio_streaming_source_data,  --                       .data
			avalon_streaming_source_valid => output_switcher_1_audio_streaming_source_valid  --                       .valid
		);

	spi_system_0 : component SPI_System
		port map (
			clk                => pll_0_outclk0_clk,                                     --         clock.clk
			reset_n            => rst_controller_reset_out_reset_ports_inv,              --         reset.reset_n
			AM_Addr            => spi_system_0_avalon_master_address,                    -- avalon_master.address
			AM_BurstCount      => spi_system_0_avalon_master_burstcount,                 --              .burstcount
			AM_ByteEnable      => spi_system_0_avalon_master_byteenable,                 --              .byteenable
			AM_DataWrite       => spi_system_0_avalon_master_writedata,                  --              .writedata
			AM_WaitRequest     => spi_system_0_avalon_master_waitrequest,                --              .waitrequest
			AM_Write           => spi_system_0_avalon_master_write,                      --              .write
			AS_Write           => mm_interconnect_1_spi_system_0_avalon_slave_write,     --  avalon_slave.write
			AS_Read            => mm_interconnect_1_spi_system_0_avalon_slave_read,      --              .read
			AS_ReadData        => mm_interconnect_1_spi_system_0_avalon_slave_readdata,  --              .readdata
			AS_WriteData       => mm_interconnect_1_spi_system_0_avalon_slave_writedata, --              .writedata
			AS_Addr            => mm_interconnect_1_spi_system_0_avalon_slave_address,   --              .address
			CONVST0            => spi_system_0_spi_interface_convst0,                    -- spi_interface.convst0
			CONVST1            => spi_system_0_spi_interface_convst1,                    --              .convst1
			CONVST2            => spi_system_0_spi_interface_convst2,                    --              .convst2
			CS0_n              => spi_system_0_spi_interface_cs0_n,                      --              .cs0_n
			CS1_n              => spi_system_0_spi_interface_cs1_n,                      --              .cs1_n
			CS2_n              => spi_system_0_spi_interface_cs2_n,                      --              .cs2_n
			MISO_00            => spi_system_0_spi_interface_miso_00,                    --              .miso_00
			MISO_01            => spi_system_0_spi_interface_miso_01,                    --              .miso_01
			MISO_10            => spi_system_0_spi_interface_miso_10,                    --              .miso_10
			MISO_11            => spi_system_0_spi_interface_miso_11,                    --              .miso_11
			MISO_20            => spi_system_0_spi_interface_miso_20,                    --              .miso_20
			MISO_21            => spi_system_0_spi_interface_miso_21,                    --              .miso_21
			Reset0             => spi_system_0_spi_interface_reset0,                     --              .reset0
			Reset1             => spi_system_0_spi_interface_reset1,                     --              .reset1
			Reset2             => spi_system_0_spi_interface_reset2,                     --              .reset2
			SCLK0              => spi_system_0_spi_interface_sclk0,                      --              .sclk0
			SCLK1              => spi_system_0_spi_interface_sclk1,                      --              .sclk1
			SCLK2              => spi_system_0_spi_interface_sclk2,                      --              .sclk2
			busy_OR0           => spi_system_0_spi_interface_busy_or0,                   --              .busy_or0
			busy_OR1           => spi_system_0_spi_interface_busy_or1,                   --              .busy_or1
			busy_OR2           => spi_system_0_spi_interface_busy_or2,                   --              .busy_or2
			Source_Data_Left   => spi_system_0_source_left_data,                         --   Source_Left.data
			Source_sop_Left    => spi_system_0_source_left_startofpacket,                --              .startofpacket
			Source_eop_Left    => spi_system_0_source_left_endofpacket,                  --              .endofpacket
			Source_Valid_Left  => spi_system_0_source_left_valid,                        --              .valid
			Source_Ready_Left  => spi_system_0_source_left_ready,                        --              .ready
			Source_Data_Right  => spi_system_0_source_right_data,                        --  Source_Right.data
			Source_Ready_Right => spi_system_0_source_right_ready,                       --              .ready
			Source_Valid_Right => spi_system_0_source_right_valid,                       --              .valid
			Source_eop_Right   => spi_system_0_source_right_endofpacket,                 --              .endofpacket
			Source_sop_Right   => spi_system_0_source_right_startofpacket                --              .startofpacket
		);

	audio_and_video_config_0 : component Pyramic_Array_audio_and_video_config_0
		port map (
			clk         => pll_0_outclk0_clk,                                                             --                    clk.clk
			reset       => rst_controller_reset_out_reset,                                                --                  reset.reset
			address     => mm_interconnect_1_audio_and_video_config_0_avalon_av_config_slave_address,     -- avalon_av_config_slave.address
			byteenable  => mm_interconnect_1_audio_and_video_config_0_avalon_av_config_slave_byteenable,  --                       .byteenable
			read        => mm_interconnect_1_audio_and_video_config_0_avalon_av_config_slave_read,        --                       .read
			write       => mm_interconnect_1_audio_and_video_config_0_avalon_av_config_slave_write,       --                       .write
			writedata   => mm_interconnect_1_audio_and_video_config_0_avalon_av_config_slave_writedata,   --                       .writedata
			readdata    => mm_interconnect_1_audio_and_video_config_0_avalon_av_config_slave_readdata,    --                       .readdata
			waitrequest => mm_interconnect_1_audio_and_video_config_0_avalon_av_config_slave_waitrequest, --                       .waitrequest
			I2C_SDAT    => audio_and_video_config_0_external_interface_SDAT,                              --     external_interface.export
			I2C_SCLK    => audio_and_video_config_0_external_interface_SCLK                               --                       .export
		);

	audio_controller : component Pyramic_Array_audio_controller
		port map (
			clk                          => pll_0_outclk0_clk,                              --                         clk.clk
			reset                        => rst_controller_reset_out_reset,                 --                       reset.reset
			from_adc_left_channel_ready  => open,                                           --  avalon_left_channel_source.ready
			from_adc_left_channel_data   => open,                                           --                            .data
			from_adc_left_channel_valid  => open,                                           --                            .valid
			from_adc_right_channel_ready => open,                                           -- avalon_right_channel_source.ready
			from_adc_right_channel_data  => open,                                           --                            .data
			from_adc_right_channel_valid => open,                                           --                            .valid
			to_dac_left_channel_data     => output_switcher_0_audio_streaming_source_data,  --    avalon_left_channel_sink.data
			to_dac_left_channel_valid    => output_switcher_0_audio_streaming_source_valid, --                            .valid
			to_dac_left_channel_ready    => output_switcher_0_audio_streaming_source_ready, --                            .ready
			to_dac_right_channel_data    => output_switcher_1_audio_streaming_source_data,  --   avalon_right_channel_sink.data
			to_dac_right_channel_valid   => output_switcher_1_audio_streaming_source_valid, --                            .valid
			to_dac_right_channel_ready   => output_switcher_1_audio_streaming_source_ready, --                            .ready
			AUD_BCLK                     => audio_0_external_interface_BCLK,                --          external_interface.export
			AUD_DACDAT                   => audio_0_external_interface_DACDAT,              --                            .export
			AUD_DACLRCK                  => audio_0_external_interface_DACLRCK              --                            .export
		);

	hps_0 : component Pyramic_Array_hps_0
		generic map (
			F2S_Width => 0,
			S2F_Width => 0
		)
		port map (
			mem_a                    => hps_0_ddr_mem_a,                                       --            memory.mem_a
			mem_ba                   => hps_0_ddr_mem_ba,                                      --                  .mem_ba
			mem_ck                   => hps_0_ddr_mem_ck,                                      --                  .mem_ck
			mem_ck_n                 => hps_0_ddr_mem_ck_n,                                    --                  .mem_ck_n
			mem_cke                  => hps_0_ddr_mem_cke,                                     --                  .mem_cke
			mem_cs_n                 => hps_0_ddr_mem_cs_n,                                    --                  .mem_cs_n
			mem_ras_n                => hps_0_ddr_mem_ras_n,                                   --                  .mem_ras_n
			mem_cas_n                => hps_0_ddr_mem_cas_n,                                   --                  .mem_cas_n
			mem_we_n                 => hps_0_ddr_mem_we_n,                                    --                  .mem_we_n
			mem_reset_n              => hps_0_ddr_mem_reset_n,                                 --                  .mem_reset_n
			mem_dq                   => hps_0_ddr_mem_dq,                                      --                  .mem_dq
			mem_dqs                  => hps_0_ddr_mem_dqs,                                     --                  .mem_dqs
			mem_dqs_n                => hps_0_ddr_mem_dqs_n,                                   --                  .mem_dqs_n
			mem_odt                  => hps_0_ddr_mem_odt,                                     --                  .mem_odt
			mem_dm                   => hps_0_ddr_mem_dm,                                      --                  .mem_dm
			oct_rzqin                => hps_0_ddr_oct_rzqin,                                   --                  .oct_rzqin
			hps_io_emac1_inst_TX_CLK => hps_0_io_hps_io_emac1_inst_TX_CLK,                     --            hps_io.hps_io_emac1_inst_TX_CLK
			hps_io_emac1_inst_TXD0   => hps_0_io_hps_io_emac1_inst_TXD0,                       --                  .hps_io_emac1_inst_TXD0
			hps_io_emac1_inst_TXD1   => hps_0_io_hps_io_emac1_inst_TXD1,                       --                  .hps_io_emac1_inst_TXD1
			hps_io_emac1_inst_TXD2   => hps_0_io_hps_io_emac1_inst_TXD2,                       --                  .hps_io_emac1_inst_TXD2
			hps_io_emac1_inst_TXD3   => hps_0_io_hps_io_emac1_inst_TXD3,                       --                  .hps_io_emac1_inst_TXD3
			hps_io_emac1_inst_RXD0   => hps_0_io_hps_io_emac1_inst_RXD0,                       --                  .hps_io_emac1_inst_RXD0
			hps_io_emac1_inst_MDIO   => hps_0_io_hps_io_emac1_inst_MDIO,                       --                  .hps_io_emac1_inst_MDIO
			hps_io_emac1_inst_MDC    => hps_0_io_hps_io_emac1_inst_MDC,                        --                  .hps_io_emac1_inst_MDC
			hps_io_emac1_inst_RX_CTL => hps_0_io_hps_io_emac1_inst_RX_CTL,                     --                  .hps_io_emac1_inst_RX_CTL
			hps_io_emac1_inst_TX_CTL => hps_0_io_hps_io_emac1_inst_TX_CTL,                     --                  .hps_io_emac1_inst_TX_CTL
			hps_io_emac1_inst_RX_CLK => hps_0_io_hps_io_emac1_inst_RX_CLK,                     --                  .hps_io_emac1_inst_RX_CLK
			hps_io_emac1_inst_RXD1   => hps_0_io_hps_io_emac1_inst_RXD1,                       --                  .hps_io_emac1_inst_RXD1
			hps_io_emac1_inst_RXD2   => hps_0_io_hps_io_emac1_inst_RXD2,                       --                  .hps_io_emac1_inst_RXD2
			hps_io_emac1_inst_RXD3   => hps_0_io_hps_io_emac1_inst_RXD3,                       --                  .hps_io_emac1_inst_RXD3
			hps_io_sdio_inst_CMD     => hps_0_io_hps_io_sdio_inst_CMD,                         --                  .hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0      => hps_0_io_hps_io_sdio_inst_D0,                          --                  .hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1      => hps_0_io_hps_io_sdio_inst_D1,                          --                  .hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK     => hps_0_io_hps_io_sdio_inst_CLK,                         --                  .hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2      => hps_0_io_hps_io_sdio_inst_D2,                          --                  .hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3      => hps_0_io_hps_io_sdio_inst_D3,                          --                  .hps_io_sdio_inst_D3
			hps_io_uart0_inst_RX     => hps_0_io_hps_io_uart0_inst_RX,                         --                  .hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX     => hps_0_io_hps_io_uart0_inst_TX,                         --                  .hps_io_uart0_inst_TX
			hps_io_gpio_inst_GPIO35  => hps_0_io_hps_io_gpio_inst_GPIO35,                      --                  .hps_io_gpio_inst_GPIO35
			hps_io_gpio_inst_GPIO53  => hps_0_io_hps_io_gpio_inst_GPIO53,                      --                  .hps_io_gpio_inst_GPIO53
			hps_io_gpio_inst_GPIO54  => hps_0_io_hps_io_gpio_inst_GPIO54,                      --                  .hps_io_gpio_inst_GPIO54
			h2f_rst_n                => hps_0_h2f_reset_reset,                                 --         h2f_reset.reset_n
			f2h_sdram0_clk           => pll_0_outclk0_clk,                                     --  f2h_sdram0_clock.clk
			f2h_sdram0_ADDRESS       => mm_interconnect_0_hps_0_f2h_sdram0_data_address,       --   f2h_sdram0_data.address
			f2h_sdram0_BURSTCOUNT    => mm_interconnect_0_hps_0_f2h_sdram0_data_burstcount,    --                  .burstcount
			f2h_sdram0_WAITREQUEST   => mm_interconnect_0_hps_0_f2h_sdram0_data_waitrequest,   --                  .waitrequest
			f2h_sdram0_READDATA      => mm_interconnect_0_hps_0_f2h_sdram0_data_readdata,      --                  .readdata
			f2h_sdram0_READDATAVALID => mm_interconnect_0_hps_0_f2h_sdram0_data_readdatavalid, --                  .readdatavalid
			f2h_sdram0_READ          => mm_interconnect_0_hps_0_f2h_sdram0_data_read,          --                  .read
			f2h_sdram0_WRITEDATA     => mm_interconnect_0_hps_0_f2h_sdram0_data_writedata,     --                  .writedata
			f2h_sdram0_BYTEENABLE    => mm_interconnect_0_hps_0_f2h_sdram0_data_byteenable,    --                  .byteenable
			f2h_sdram0_WRITE         => mm_interconnect_0_hps_0_f2h_sdram0_data_write,         --                  .write
			h2f_lw_axi_clk           => pll_0_outclk0_clk,                                     --  h2f_lw_axi_clock.clk
			h2f_lw_AWID              => hps_0_h2f_lw_axi_master_awid,                          -- h2f_lw_axi_master.awid
			h2f_lw_AWADDR            => hps_0_h2f_lw_axi_master_awaddr,                        --                  .awaddr
			h2f_lw_AWLEN             => hps_0_h2f_lw_axi_master_awlen,                         --                  .awlen
			h2f_lw_AWSIZE            => hps_0_h2f_lw_axi_master_awsize,                        --                  .awsize
			h2f_lw_AWBURST           => hps_0_h2f_lw_axi_master_awburst,                       --                  .awburst
			h2f_lw_AWLOCK            => hps_0_h2f_lw_axi_master_awlock,                        --                  .awlock
			h2f_lw_AWCACHE           => hps_0_h2f_lw_axi_master_awcache,                       --                  .awcache
			h2f_lw_AWPROT            => hps_0_h2f_lw_axi_master_awprot,                        --                  .awprot
			h2f_lw_AWVALID           => hps_0_h2f_lw_axi_master_awvalid,                       --                  .awvalid
			h2f_lw_AWREADY           => hps_0_h2f_lw_axi_master_awready,                       --                  .awready
			h2f_lw_WID               => hps_0_h2f_lw_axi_master_wid,                           --                  .wid
			h2f_lw_WDATA             => hps_0_h2f_lw_axi_master_wdata,                         --                  .wdata
			h2f_lw_WSTRB             => hps_0_h2f_lw_axi_master_wstrb,                         --                  .wstrb
			h2f_lw_WLAST             => hps_0_h2f_lw_axi_master_wlast,                         --                  .wlast
			h2f_lw_WVALID            => hps_0_h2f_lw_axi_master_wvalid,                        --                  .wvalid
			h2f_lw_WREADY            => hps_0_h2f_lw_axi_master_wready,                        --                  .wready
			h2f_lw_BID               => hps_0_h2f_lw_axi_master_bid,                           --                  .bid
			h2f_lw_BRESP             => hps_0_h2f_lw_axi_master_bresp,                         --                  .bresp
			h2f_lw_BVALID            => hps_0_h2f_lw_axi_master_bvalid,                        --                  .bvalid
			h2f_lw_BREADY            => hps_0_h2f_lw_axi_master_bready,                        --                  .bready
			h2f_lw_ARID              => hps_0_h2f_lw_axi_master_arid,                          --                  .arid
			h2f_lw_ARADDR            => hps_0_h2f_lw_axi_master_araddr,                        --                  .araddr
			h2f_lw_ARLEN             => hps_0_h2f_lw_axi_master_arlen,                         --                  .arlen
			h2f_lw_ARSIZE            => hps_0_h2f_lw_axi_master_arsize,                        --                  .arsize
			h2f_lw_ARBURST           => hps_0_h2f_lw_axi_master_arburst,                       --                  .arburst
			h2f_lw_ARLOCK            => hps_0_h2f_lw_axi_master_arlock,                        --                  .arlock
			h2f_lw_ARCACHE           => hps_0_h2f_lw_axi_master_arcache,                       --                  .arcache
			h2f_lw_ARPROT            => hps_0_h2f_lw_axi_master_arprot,                        --                  .arprot
			h2f_lw_ARVALID           => hps_0_h2f_lw_axi_master_arvalid,                       --                  .arvalid
			h2f_lw_ARREADY           => hps_0_h2f_lw_axi_master_arready,                       --                  .arready
			h2f_lw_RID               => hps_0_h2f_lw_axi_master_rid,                           --                  .rid
			h2f_lw_RDATA             => hps_0_h2f_lw_axi_master_rdata,                         --                  .rdata
			h2f_lw_RRESP             => hps_0_h2f_lw_axi_master_rresp,                         --                  .rresp
			h2f_lw_RLAST             => hps_0_h2f_lw_axi_master_rlast,                         --                  .rlast
			h2f_lw_RVALID            => hps_0_h2f_lw_axi_master_rvalid,                        --                  .rvalid
			h2f_lw_RREADY            => hps_0_h2f_lw_axi_master_rready                         --                  .rready
		);

	jtag_uart_0 : component Pyramic_Array_jtag_uart_0
		port map (
			clk            => pll_0_outclk0_clk,                            --               clk.clk
			rst_n          => rst_controller_001_reset_out_reset_ports_inv, --             reset.reset_n
			av_chipselect  => open,                                         -- avalon_jtag_slave.chipselect
			av_address     => open,                                         --                  .address
			av_read_n      => open,                                         --                  .read_n
			av_readdata    => open,                                         --                  .readdata
			av_write_n     => open,                                         --                  .write_n
			av_writedata   => open,                                         --                  .writedata
			av_waitrequest => open,                                         --                  .waitrequest
			av_irq         => open                                          --               irq.irq
		);

	pll_0 : component Pyramic_Array_pll_0
		port map (
			refclk   => clk_clk,                            --  refclk.clk
			rst      => rst_controller_002_reset_out_reset, --   reset.reset
			outclk_0 => pll_0_outclk0_clk,                  -- outclk0.clk
			outclk_1 => open,                               -- outclk1.clk
			outclk_2 => pll_0_sdram_clk,                    -- outclk2.clk
			outclk_3 => open,                               -- outclk3.clk
			locked   => open                                -- (terminated)
		);

	pll_1 : component Pyramic_Array_pll_1
		port map (
			refclk   => pll_0_outclk0_clk,       --  refclk.clk
			rst      => reset_reset_n_ports_inv, --   reset.reset
			outclk_0 => pll_0_outclk3_audio_clk, -- outclk0.clk
			locked   => open                     --  locked.export
		);

	sysid : component Pyramic_Array_sysid
		port map (
			clock    => pll_0_outclk0_clk,                            --           clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv, --         reset.reset_n
			readdata => open,                                         -- control_slave.readdata
			address  => open                                          --              .address
		);

	mm_interconnect_0 : component Pyramic_Array_mm_interconnect_0
		port map (
			pll_0_outclk0_clk                                                  => pll_0_outclk0_clk,                                     --                                                pll_0_outclk0.clk
			hps_0_f2h_sdram0_data_translator_reset_reset_bridge_in_reset_reset => rst_controller_003_reset_out_reset,                    -- hps_0_f2h_sdram0_data_translator_reset_reset_bridge_in_reset.reset
			Output_Switcher_0_reset_reset_bridge_in_reset_reset                => rst_controller_reset_out_reset,                        --                Output_Switcher_0_reset_reset_bridge_in_reset.reset
			Output_Switcher_0_DMA_address                                      => output_switcher_0_dma_address,                         --                                        Output_Switcher_0_DMA.address
			Output_Switcher_0_DMA_waitrequest                                  => output_switcher_0_dma_waitrequest,                     --                                                             .waitrequest
			Output_Switcher_0_DMA_byteenable                                   => output_switcher_0_dma_byteenable,                      --                                                             .byteenable
			Output_Switcher_0_DMA_read                                         => output_switcher_0_dma_read,                            --                                                             .read
			Output_Switcher_0_DMA_readdata                                     => output_switcher_0_dma_readdata,                        --                                                             .readdata
			Output_Switcher_0_DMA_readdatavalid                                => output_switcher_0_dma_readdatavalid,                   --                                                             .readdatavalid
			Output_Switcher_1_DMA_address                                      => output_switcher_1_dma_address,                         --                                        Output_Switcher_1_DMA.address
			Output_Switcher_1_DMA_waitrequest                                  => output_switcher_1_dma_waitrequest,                     --                                                             .waitrequest
			Output_Switcher_1_DMA_byteenable                                   => output_switcher_1_dma_byteenable,                      --                                                             .byteenable
			Output_Switcher_1_DMA_read                                         => output_switcher_1_dma_read,                            --                                                             .read
			Output_Switcher_1_DMA_readdata                                     => output_switcher_1_dma_readdata,                        --                                                             .readdata
			Output_Switcher_1_DMA_readdatavalid                                => output_switcher_1_dma_readdatavalid,                   --                                                             .readdatavalid
			SPI_System_0_avalon_master_address                                 => spi_system_0_avalon_master_address,                    --                                   SPI_System_0_avalon_master.address
			SPI_System_0_avalon_master_waitrequest                             => spi_system_0_avalon_master_waitrequest,                --                                                             .waitrequest
			SPI_System_0_avalon_master_burstcount                              => spi_system_0_avalon_master_burstcount,                 --                                                             .burstcount
			SPI_System_0_avalon_master_byteenable                              => spi_system_0_avalon_master_byteenable,                 --                                                             .byteenable
			SPI_System_0_avalon_master_write                                   => spi_system_0_avalon_master_write,                      --                                                             .write
			SPI_System_0_avalon_master_writedata                               => spi_system_0_avalon_master_writedata,                  --                                                             .writedata
			hps_0_f2h_sdram0_data_address                                      => mm_interconnect_0_hps_0_f2h_sdram0_data_address,       --                                        hps_0_f2h_sdram0_data.address
			hps_0_f2h_sdram0_data_write                                        => mm_interconnect_0_hps_0_f2h_sdram0_data_write,         --                                                             .write
			hps_0_f2h_sdram0_data_read                                         => mm_interconnect_0_hps_0_f2h_sdram0_data_read,          --                                                             .read
			hps_0_f2h_sdram0_data_readdata                                     => mm_interconnect_0_hps_0_f2h_sdram0_data_readdata,      --                                                             .readdata
			hps_0_f2h_sdram0_data_writedata                                    => mm_interconnect_0_hps_0_f2h_sdram0_data_writedata,     --                                                             .writedata
			hps_0_f2h_sdram0_data_burstcount                                   => mm_interconnect_0_hps_0_f2h_sdram0_data_burstcount,    --                                                             .burstcount
			hps_0_f2h_sdram0_data_byteenable                                   => mm_interconnect_0_hps_0_f2h_sdram0_data_byteenable,    --                                                             .byteenable
			hps_0_f2h_sdram0_data_readdatavalid                                => mm_interconnect_0_hps_0_f2h_sdram0_data_readdatavalid, --                                                             .readdatavalid
			hps_0_f2h_sdram0_data_waitrequest                                  => mm_interconnect_0_hps_0_f2h_sdram0_data_waitrequest    --                                                             .waitrequest
		);

	mm_interconnect_1 : component Pyramic_Array_mm_interconnect_1
		port map (
			hps_0_h2f_lw_axi_master_awid                                        => hps_0_h2f_lw_axi_master_awid,                                                  --                                       hps_0_h2f_lw_axi_master.awid
			hps_0_h2f_lw_axi_master_awaddr                                      => hps_0_h2f_lw_axi_master_awaddr,                                                --                                                              .awaddr
			hps_0_h2f_lw_axi_master_awlen                                       => hps_0_h2f_lw_axi_master_awlen,                                                 --                                                              .awlen
			hps_0_h2f_lw_axi_master_awsize                                      => hps_0_h2f_lw_axi_master_awsize,                                                --                                                              .awsize
			hps_0_h2f_lw_axi_master_awburst                                     => hps_0_h2f_lw_axi_master_awburst,                                               --                                                              .awburst
			hps_0_h2f_lw_axi_master_awlock                                      => hps_0_h2f_lw_axi_master_awlock,                                                --                                                              .awlock
			hps_0_h2f_lw_axi_master_awcache                                     => hps_0_h2f_lw_axi_master_awcache,                                               --                                                              .awcache
			hps_0_h2f_lw_axi_master_awprot                                      => hps_0_h2f_lw_axi_master_awprot,                                                --                                                              .awprot
			hps_0_h2f_lw_axi_master_awvalid                                     => hps_0_h2f_lw_axi_master_awvalid,                                               --                                                              .awvalid
			hps_0_h2f_lw_axi_master_awready                                     => hps_0_h2f_lw_axi_master_awready,                                               --                                                              .awready
			hps_0_h2f_lw_axi_master_wid                                         => hps_0_h2f_lw_axi_master_wid,                                                   --                                                              .wid
			hps_0_h2f_lw_axi_master_wdata                                       => hps_0_h2f_lw_axi_master_wdata,                                                 --                                                              .wdata
			hps_0_h2f_lw_axi_master_wstrb                                       => hps_0_h2f_lw_axi_master_wstrb,                                                 --                                                              .wstrb
			hps_0_h2f_lw_axi_master_wlast                                       => hps_0_h2f_lw_axi_master_wlast,                                                 --                                                              .wlast
			hps_0_h2f_lw_axi_master_wvalid                                      => hps_0_h2f_lw_axi_master_wvalid,                                                --                                                              .wvalid
			hps_0_h2f_lw_axi_master_wready                                      => hps_0_h2f_lw_axi_master_wready,                                                --                                                              .wready
			hps_0_h2f_lw_axi_master_bid                                         => hps_0_h2f_lw_axi_master_bid,                                                   --                                                              .bid
			hps_0_h2f_lw_axi_master_bresp                                       => hps_0_h2f_lw_axi_master_bresp,                                                 --                                                              .bresp
			hps_0_h2f_lw_axi_master_bvalid                                      => hps_0_h2f_lw_axi_master_bvalid,                                                --                                                              .bvalid
			hps_0_h2f_lw_axi_master_bready                                      => hps_0_h2f_lw_axi_master_bready,                                                --                                                              .bready
			hps_0_h2f_lw_axi_master_arid                                        => hps_0_h2f_lw_axi_master_arid,                                                  --                                                              .arid
			hps_0_h2f_lw_axi_master_araddr                                      => hps_0_h2f_lw_axi_master_araddr,                                                --                                                              .araddr
			hps_0_h2f_lw_axi_master_arlen                                       => hps_0_h2f_lw_axi_master_arlen,                                                 --                                                              .arlen
			hps_0_h2f_lw_axi_master_arsize                                      => hps_0_h2f_lw_axi_master_arsize,                                                --                                                              .arsize
			hps_0_h2f_lw_axi_master_arburst                                     => hps_0_h2f_lw_axi_master_arburst,                                               --                                                              .arburst
			hps_0_h2f_lw_axi_master_arlock                                      => hps_0_h2f_lw_axi_master_arlock,                                                --                                                              .arlock
			hps_0_h2f_lw_axi_master_arcache                                     => hps_0_h2f_lw_axi_master_arcache,                                               --                                                              .arcache
			hps_0_h2f_lw_axi_master_arprot                                      => hps_0_h2f_lw_axi_master_arprot,                                                --                                                              .arprot
			hps_0_h2f_lw_axi_master_arvalid                                     => hps_0_h2f_lw_axi_master_arvalid,                                               --                                                              .arvalid
			hps_0_h2f_lw_axi_master_arready                                     => hps_0_h2f_lw_axi_master_arready,                                               --                                                              .arready
			hps_0_h2f_lw_axi_master_rid                                         => hps_0_h2f_lw_axi_master_rid,                                                   --                                                              .rid
			hps_0_h2f_lw_axi_master_rdata                                       => hps_0_h2f_lw_axi_master_rdata,                                                 --                                                              .rdata
			hps_0_h2f_lw_axi_master_rresp                                       => hps_0_h2f_lw_axi_master_rresp,                                                 --                                                              .rresp
			hps_0_h2f_lw_axi_master_rlast                                       => hps_0_h2f_lw_axi_master_rlast,                                                 --                                                              .rlast
			hps_0_h2f_lw_axi_master_rvalid                                      => hps_0_h2f_lw_axi_master_rvalid,                                                --                                                              .rvalid
			hps_0_h2f_lw_axi_master_rready                                      => hps_0_h2f_lw_axi_master_rready,                                                --                                                              .rready
			pll_0_outclk0_clk                                                   => pll_0_outclk0_clk,                                                             --                                                 pll_0_outclk0.clk
			audio_and_video_config_0_reset_reset_bridge_in_reset_reset          => rst_controller_reset_out_reset,                                                --          audio_and_video_config_0_reset_reset_bridge_in_reset.reset
			hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset => rst_controller_003_reset_out_reset,                                            -- hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
			audio_and_video_config_0_avalon_av_config_slave_address             => mm_interconnect_1_audio_and_video_config_0_avalon_av_config_slave_address,     --               audio_and_video_config_0_avalon_av_config_slave.address
			audio_and_video_config_0_avalon_av_config_slave_write               => mm_interconnect_1_audio_and_video_config_0_avalon_av_config_slave_write,       --                                                              .write
			audio_and_video_config_0_avalon_av_config_slave_read                => mm_interconnect_1_audio_and_video_config_0_avalon_av_config_slave_read,        --                                                              .read
			audio_and_video_config_0_avalon_av_config_slave_readdata            => mm_interconnect_1_audio_and_video_config_0_avalon_av_config_slave_readdata,    --                                                              .readdata
			audio_and_video_config_0_avalon_av_config_slave_writedata           => mm_interconnect_1_audio_and_video_config_0_avalon_av_config_slave_writedata,   --                                                              .writedata
			audio_and_video_config_0_avalon_av_config_slave_byteenable          => mm_interconnect_1_audio_and_video_config_0_avalon_av_config_slave_byteenable,  --                                                              .byteenable
			audio_and_video_config_0_avalon_av_config_slave_waitrequest         => mm_interconnect_1_audio_and_video_config_0_avalon_av_config_slave_waitrequest, --                                                              .waitrequest
			SPI_System_0_avalon_slave_address                                   => mm_interconnect_1_spi_system_0_avalon_slave_address,                           --                                     SPI_System_0_avalon_slave.address
			SPI_System_0_avalon_slave_write                                     => mm_interconnect_1_spi_system_0_avalon_slave_write,                             --                                                              .write
			SPI_System_0_avalon_slave_read                                      => mm_interconnect_1_spi_system_0_avalon_slave_read,                              --                                                              .read
			SPI_System_0_avalon_slave_readdata                                  => mm_interconnect_1_spi_system_0_avalon_slave_readdata,                          --                                                              .readdata
			SPI_System_0_avalon_slave_writedata                                 => mm_interconnect_1_spi_system_0_avalon_slave_writedata                          --                                                              .writedata
		);

	avalon_st_adapter : component Pyramic_Array_avalon_st_adapter
		generic map (
			inBitsPerSymbol => 22,
			inUsePackets    => 1,
			inDataWidth     => 22,
			inChannelWidth  => 0,
			inErrorWidth    => 0,
			inUseEmptyPort  => 0,
			inUseValid      => 1,
			inUseReady      => 1,
			inReadyLatency  => 0,
			outDataWidth    => 22,
			outChannelWidth => 0,
			outErrorWidth   => 2,
			outUseEmptyPort => 0,
			outUseValid     => 1,
			outUseReady     => 0,
			outReadyLatency => 0
		)
		port map (
			in_clk_0_clk        => pll_0_outclk0_clk,                      -- in_clk_0.clk
			in_rst_0_reset      => rst_controller_reset_out_reset,         -- in_rst_0.reset
			in_0_data           => spi_system_0_source_left_data,          --     in_0.data
			in_0_valid          => spi_system_0_source_left_valid,         --         .valid
			in_0_ready          => spi_system_0_source_left_ready,         --         .ready
			in_0_startofpacket  => spi_system_0_source_left_startofpacket, --         .startofpacket
			in_0_endofpacket    => spi_system_0_source_left_endofpacket,   --         .endofpacket
			out_0_data          => avalon_st_adapter_out_0_data,           --    out_0.data
			out_0_valid         => avalon_st_adapter_out_0_valid,          --         .valid
			out_0_startofpacket => avalon_st_adapter_out_0_startofpacket,  --         .startofpacket
			out_0_endofpacket   => avalon_st_adapter_out_0_endofpacket,    --         .endofpacket
			out_0_error         => avalon_st_adapter_out_0_error           --         .error
		);

	avalon_st_adapter_001 : component Pyramic_Array_avalon_st_adapter
		generic map (
			inBitsPerSymbol => 22,
			inUsePackets    => 1,
			inDataWidth     => 22,
			inChannelWidth  => 0,
			inErrorWidth    => 0,
			inUseEmptyPort  => 0,
			inUseValid      => 1,
			inUseReady      => 1,
			inReadyLatency  => 0,
			outDataWidth    => 22,
			outChannelWidth => 0,
			outErrorWidth   => 2,
			outUseEmptyPort => 0,
			outUseValid     => 1,
			outUseReady     => 0,
			outReadyLatency => 0
		)
		port map (
			in_clk_0_clk        => pll_0_outclk0_clk,                         -- in_clk_0.clk
			in_rst_0_reset      => rst_controller_reset_out_reset,            -- in_rst_0.reset
			in_0_data           => spi_system_0_source_right_data,            --     in_0.data
			in_0_valid          => spi_system_0_source_right_valid,           --         .valid
			in_0_ready          => spi_system_0_source_right_ready,           --         .ready
			in_0_startofpacket  => spi_system_0_source_right_startofpacket,   --         .startofpacket
			in_0_endofpacket    => spi_system_0_source_right_endofpacket,     --         .endofpacket
			out_0_data          => avalon_st_adapter_001_out_0_data,          --    out_0.data
			out_0_valid         => avalon_st_adapter_001_out_0_valid,         --         .valid
			out_0_startofpacket => avalon_st_adapter_001_out_0_startofpacket, --         .startofpacket
			out_0_endofpacket   => avalon_st_adapter_001_out_0_endofpacket,   --         .endofpacket
			out_0_error         => avalon_st_adapter_001_out_0_error          --         .error
		);

	avalon_st_adapter_002 : component Pyramic_Array_avalon_st_adapter_002
		generic map (
			inBitsPerSymbol => 32,
			inUsePackets    => 1,
			inDataWidth     => 32,
			inChannelWidth  => 6,
			inErrorWidth    => 2,
			inUseEmptyPort  => 0,
			inUseValid      => 1,
			inUseReady      => 0,
			inReadyLatency  => 0,
			outDataWidth    => 32,
			outChannelWidth => 6,
			outErrorWidth   => 0,
			outUseEmptyPort => 0,
			outUseValid     => 1,
			outUseReady     => 1,
			outReadyLatency => 0
		)
		port map (
			in_clk_0_clk        => pll_0_outclk0_clk,                              -- in_clk_0.clk
			in_rst_0_reset      => rst_controller_reset_out_reset,                 -- in_rst_0.reset
			in_0_data           => fir_left_avalon_streaming_source_data,          --     in_0.data
			in_0_valid          => fir_left_avalon_streaming_source_valid,         --         .valid
			in_0_startofpacket  => fir_left_avalon_streaming_source_startofpacket, --         .startofpacket
			in_0_endofpacket    => fir_left_avalon_streaming_source_endofpacket,   --         .endofpacket
			in_0_error          => fir_left_avalon_streaming_source_error,         --         .error
			in_0_channel        => fir_left_avalon_streaming_source_channel,       --         .channel
			out_0_data          => avalon_st_adapter_002_out_0_data,               --    out_0.data
			out_0_valid         => avalon_st_adapter_002_out_0_valid,              --         .valid
			out_0_ready         => avalon_st_adapter_002_out_0_ready,              --         .ready
			out_0_startofpacket => avalon_st_adapter_002_out_0_startofpacket,      --         .startofpacket
			out_0_endofpacket   => avalon_st_adapter_002_out_0_endofpacket,        --         .endofpacket
			out_0_channel       => avalon_st_adapter_002_out_0_channel             --         .channel
		);

	avalon_st_adapter_003 : component Pyramic_Array_avalon_st_adapter_002
		generic map (
			inBitsPerSymbol => 32,
			inUsePackets    => 1,
			inDataWidth     => 32,
			inChannelWidth  => 6,
			inErrorWidth    => 2,
			inUseEmptyPort  => 0,
			inUseValid      => 1,
			inUseReady      => 0,
			inReadyLatency  => 0,
			outDataWidth    => 32,
			outChannelWidth => 6,
			outErrorWidth   => 0,
			outUseEmptyPort => 0,
			outUseValid     => 1,
			outUseReady     => 1,
			outReadyLatency => 0
		)
		port map (
			in_clk_0_clk        => pll_0_outclk0_clk,                               -- in_clk_0.clk
			in_rst_0_reset      => rst_controller_reset_out_reset,                  -- in_rst_0.reset
			in_0_data           => fir_right_avalon_streaming_source_data,          --     in_0.data
			in_0_valid          => fir_right_avalon_streaming_source_valid,         --         .valid
			in_0_startofpacket  => fir_right_avalon_streaming_source_startofpacket, --         .startofpacket
			in_0_endofpacket    => fir_right_avalon_streaming_source_endofpacket,   --         .endofpacket
			in_0_error          => fir_right_avalon_streaming_source_error,         --         .error
			in_0_channel        => fir_right_avalon_streaming_source_channel,       --         .channel
			out_0_data          => avalon_st_adapter_003_out_0_data,                --    out_0.data
			out_0_valid         => avalon_st_adapter_003_out_0_valid,               --         .valid
			out_0_ready         => avalon_st_adapter_003_out_0_ready,               --         .ready
			out_0_startofpacket => avalon_st_adapter_003_out_0_startofpacket,       --         .startofpacket
			out_0_endofpacket   => avalon_st_adapter_003_out_0_endofpacket,         --         .endofpacket
			out_0_channel       => avalon_st_adapter_003_out_0_channel              --         .channel
		);

	rst_controller : component pyramic_array_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => pll_0_outclk0_clk,              --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component pyramic_array_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => hps_0_h2f_reset_reset_ports_inv,    -- reset_in1.reset
			clk            => pll_0_outclk0_clk,                  --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_002 : component pyramic_array_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "none",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => hps_0_h2f_reset_reset_ports_inv,    -- reset_in1.reset
			clk            => open,                               --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_003 : component pyramic_array_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => hps_0_h2f_reset_reset_ports_inv,    -- reset_in0.reset
			clk            => pll_0_outclk0_clk,                  --       clk.clk
			reset_out      => rst_controller_003_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

	hps_0_h2f_reset_reset_ports_inv <= not hps_0_h2f_reset_reset;

end architecture rtl; -- of Pyramic_Array
